// niosII_system.v

// Generated using ACDS version 12.1sp1 243 at 2017.03.26.17:18:02

`timescale 1 ps / 1 ps
module niosII_system (
		input  wire        reset_0_reset_n,                                                                  //                                     reset_0.reset_n
		output wire        altpll_0_c0_clk,                                                                  //                                 altpll_0_c0.clk
		output wire [0:0]  tristate_conduit_bridge_0_out_generic_tristate_controller_0_tcm_read_n_out,       //               tristate_conduit_bridge_0_out.generic_tristate_controller_0_tcm_read_n_out
		inout  wire [7:0]  tristate_conduit_bridge_0_out_generic_tristate_controller_0_tcm_data_out,         //                                            .generic_tristate_controller_0_tcm_data_out
		output wire [0:0]  tristate_conduit_bridge_0_out_generic_tristate_controller_0_tcm_chipselect_n_out, //                                            .generic_tristate_controller_0_tcm_chipselect_n_out
		output wire [0:0]  tristate_conduit_bridge_0_out_generic_tristate_controller_0_tcm_write_n_out,      //                                            .generic_tristate_controller_0_tcm_write_n_out
		output wire [21:0] tristate_conduit_bridge_0_out_generic_tristate_controller_0_tcm_address_out,      //                                            .generic_tristate_controller_0_tcm_address_out
		inout  wire        i2c_sda_external_connection_export,                                               //                 i2c_sda_external_connection.export
		inout  wire        audio_and_video_config_0_external_interface_SDAT,                                 // audio_and_video_config_0_external_interface.SDAT
		output wire        audio_and_video_config_0_external_interface_SCLK,                                 //                                            .SCLK
		input  wire        switch_external_connection_export,                                                //                  switch_external_connection.export
		input  wire        clk_clk,                                                                          //                                         clk.clk
		output wire [11:0] sdram_0_wire_addr,                                                                //                                sdram_0_wire.addr
		output wire [1:0]  sdram_0_wire_ba,                                                                  //                                            .ba
		output wire        sdram_0_wire_cas_n,                                                               //                                            .cas_n
		output wire        sdram_0_wire_cke,                                                                 //                                            .cke
		output wire        sdram_0_wire_cs_n,                                                                //                                            .cs_n
		inout  wire [15:0] sdram_0_wire_dq,                                                                  //                                            .dq
		output wire [1:0]  sdram_0_wire_dqm,                                                                 //                                            .dqm
		output wire        sdram_0_wire_ras_n,                                                               //                                            .ras_n
		output wire        sdram_0_wire_we_n,                                                                //                                            .we_n
		output wire [7:0]  green_leds_external_connection_export,                                            //              green_leds_external_connection.export
		input  wire        spi_0_external_MISO,                                                              //                              spi_0_external.MISO
		output wire        spi_0_external_MOSI,                                                              //                                            .MOSI
		output wire        spi_0_external_SCLK,                                                              //                                            .SCLK
		output wire        spi_0_external_SS_n,                                                              //                                            .SS_n
		input  wire        audio_0_external_interface_ADCDAT,                                                //                  audio_0_external_interface.ADCDAT
		input  wire        audio_0_external_interface_ADCLRCK,                                               //                                            .ADCLRCK
		input  wire        audio_0_external_interface_BCLK,                                                  //                                            .BCLK
		output wire        audio_0_external_interface_DACDAT,                                                //                                            .DACDAT
		input  wire        audio_0_external_interface_DACLRCK,                                               //                                            .DACLRCK
		output wire        i2c_scl_external_connection_export,                                               //                 i2c_scl_external_connection.export
		output wire [3:0]  drum_out_external_connection_export,                                              //                drum_out_external_connection.export
		inout  wire [7:0]  character_lcd_0_external_interface_DATA,                                          //          character_lcd_0_external_interface.DATA
		output wire        character_lcd_0_external_interface_ON,                                            //                                            .ON
		output wire        character_lcd_0_external_interface_BLON,                                          //                                            .BLON
		output wire        character_lcd_0_external_interface_EN,                                            //                                            .EN
		output wire        character_lcd_0_external_interface_RS,                                            //                                            .RS
		output wire        character_lcd_0_external_interface_RW,                                            //                                            .RW
		inout  wire        i2c_sda_2_external_connection_export,                                             //               i2c_sda_2_external_connection.export
		output wire        up_clocks_0_audio_clk_clk,                                                        //                       up_clocks_0_audio_clk.clk
		input  wire        reset_reset_n,                                                                    //                                       reset.reset_n
		input  wire        clk_1_clk,                                                                        //                                       clk_1.clk
		output wire        i2c_scl_2_external_connection_export,                                             //               i2c_scl_2_external_connection.export
		inout  wire [15:0] sram_0_external_interface_DQ,                                                     //                   sram_0_external_interface.DQ
		output wire [17:0] sram_0_external_interface_ADDR,                                                   //                                            .ADDR
		output wire        sram_0_external_interface_LB_N,                                                   //                                            .LB_N
		output wire        sram_0_external_interface_UB_N,                                                   //                                            .UB_N
		output wire        sram_0_external_interface_CE_N,                                                   //                                            .CE_N
		output wire        sram_0_external_interface_OE_N,                                                   //                                            .OE_N
		output wire        sram_0_external_interface_WE_N                                                    //                                            .WE_N
	);

	wire          altpll_0_c1_clk;                                                                                                      // altpll_0:c1 -> [I2C_SCL:clk, I2C_SCL_2:clk, I2C_SCL_2_s1_translator:clk, I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:clk, I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, I2C_SCL_s1_translator:clk, I2C_SCL_s1_translator_avalon_universal_slave_0_agent:clk, I2C_SCL_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, I2C_SDA:clk, I2C_SDA_2:clk, I2C_SDA_2_s1_translator:clk, I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:clk, I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, I2C_SDA_s1_translator:clk, I2C_SDA_s1_translator_avalon_universal_slave_0_agent:clk, I2C_SDA_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, addr_router:clk, addr_router_001:clk, burst_adapter:clk, burst_adapter_001:clk, burst_adapter_002:clk, burst_adapter_003:clk, character_lcd_0:clk, character_lcd_0_avalon_lcd_slave_translator:clk, character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:clk, character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, cmd_xbar_demux:clk, cmd_xbar_demux_001:clk, cmd_xbar_mux:clk, cmd_xbar_mux_001:clk, cmd_xbar_mux_002:clk, cmd_xbar_mux_003:clk, cmd_xbar_mux_004:clk, cmd_xbar_mux_005:clk, crosser:in_clk, crosser_001:in_clk, crosser_002:in_clk, crosser_003:out_clk, crosser_004:out_clk, crosser_005:out_clk, drum_out:clk, drum_out_s1_translator:clk, drum_out_s1_translator_avalon_universal_slave_0_agent:clk, drum_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, generic_tristate_controller_0:clk_clk, generic_tristate_controller_0_uas_translator:clk, generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:clk, generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, green_leds:clk, green_leds_s1_translator:clk, green_leds_s1_translator_avalon_universal_slave_0_agent:clk, green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, id_router:clk, id_router_001:clk, id_router_002:clk, id_router_003:clk, id_router_004:clk, id_router_005:clk, id_router_007:clk, id_router_008:clk, id_router_009:clk, id_router_010:clk, id_router_011:clk, id_router_012:clk, id_router_015:clk, id_router_016:clk, id_router_017:clk, id_router_018:clk, id_router_019:clk, irq_mapper:clk, jtag_uart_0:clk, jtag_uart_0_avalon_jtag_slave_translator:clk, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:clk, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, limiter:clk, limiter_001:clk, nios2_qsys_0:clk, nios2_qsys_0_data_master_translator:clk, nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:clk, nios2_qsys_0_instruction_master_translator:clk, nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:clk, nios2_qsys_0_jtag_debug_module_translator:clk, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:clk, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, onchip_memory2_0:clk, onchip_memory2_0_s1_translator:clk, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:clk, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rsp_xbar_demux:clk, rsp_xbar_demux_001:clk, rsp_xbar_demux_002:clk, rsp_xbar_demux_003:clk, rsp_xbar_demux_004:clk, rsp_xbar_demux_005:clk, rsp_xbar_demux_007:clk, rsp_xbar_demux_008:clk, rsp_xbar_demux_009:clk, rsp_xbar_demux_010:clk, rsp_xbar_demux_011:clk, rsp_xbar_demux_012:clk, rsp_xbar_demux_015:clk, rsp_xbar_demux_016:clk, rsp_xbar_demux_017:clk, rsp_xbar_demux_018:clk, rsp_xbar_demux_019:clk, rsp_xbar_mux:clk, rsp_xbar_mux_001:clk, rst_controller:clk, sd_card_spi_master:clk, sd_card_spi_master_spi_control_port_translator:clk, sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:clk, sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, sdram_0:clk, sdram_0_s1_translator:clk, sdram_0_s1_translator_avalon_universal_slave_0_agent:clk, sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, sram_0:clk, sram_0_avalon_sram_slave_translator:clk, sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:clk, sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, switch:clk, switch_s1_translator:clk, switch_s1_translator_avalon_universal_slave_0_agent:clk, switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, sysid_qsys_0:clock, sysid_qsys_0_control_slave_translator:clk, sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:clk, sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, timer_0:clk, timer_0_s1_translator:clk, timer_0_s1_translator_avalon_universal_slave_0_agent:clk, timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, tristate_conduit_bridge_0:clk, tristate_conduit_pin_sharer_0:clk_clk, up_clocks_0:CLOCK_50, up_clocks_1:CLOCK_50, width_adapter:clk, width_adapter_001:clk, width_adapter_002:clk, width_adapter_003:clk, width_adapter_004:clk, width_adapter_005:clk, width_adapter_006:clk, width_adapter_007:clk]
	wire          up_clocks_1_audio_clk_clk;                                                                                            // up_clocks_1:AUD_CLK -> [audio_0:clk, audio_0_avalon_audio_slave_translator:clk, audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:clk, audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, audio_and_video_config_0:clk, audio_and_video_config_0_avalon_av_config_slave_translator:clk, audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:clk, audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, crosser_001:out_clk, crosser_002:out_clk, crosser_004:in_clk, crosser_005:in_clk, id_router_013:clk, id_router_014:clk, rsp_xbar_demux_013:clk, rsp_xbar_demux_014:clk, rst_controller_002:clk]
	wire    [0:0] tristate_conduit_pin_sharer_0_tcm_generic_tristate_controller_0_tcm_read_n_out_out;                                   // tristate_conduit_pin_sharer_0:generic_tristate_controller_0_tcm_read_n_out -> tristate_conduit_bridge_0:tcs_generic_tristate_controller_0_tcm_read_n_out
	wire    [0:0] tristate_conduit_pin_sharer_0_tcm_generic_tristate_controller_0_tcm_write_n_out_out;                                  // tristate_conduit_pin_sharer_0:generic_tristate_controller_0_tcm_write_n_out -> tristate_conduit_bridge_0:tcs_generic_tristate_controller_0_tcm_write_n_out
	wire          tristate_conduit_pin_sharer_0_tcm_grant;                                                                              // tristate_conduit_bridge_0:grant -> tristate_conduit_pin_sharer_0:grant
	wire    [7:0] tristate_conduit_pin_sharer_0_tcm_generic_tristate_controller_0_tcm_data_out_in;                                      // tristate_conduit_bridge_0:tcs_generic_tristate_controller_0_tcm_data_in -> tristate_conduit_pin_sharer_0:generic_tristate_controller_0_tcm_data_in
	wire    [7:0] tristate_conduit_pin_sharer_0_tcm_generic_tristate_controller_0_tcm_data_out_out;                                     // tristate_conduit_pin_sharer_0:generic_tristate_controller_0_tcm_data_out -> tristate_conduit_bridge_0:tcs_generic_tristate_controller_0_tcm_data_out
	wire          tristate_conduit_pin_sharer_0_tcm_request;                                                                            // tristate_conduit_pin_sharer_0:request -> tristate_conduit_bridge_0:request
	wire    [0:0] tristate_conduit_pin_sharer_0_tcm_generic_tristate_controller_0_tcm_chipselect_n_out_out;                             // tristate_conduit_pin_sharer_0:generic_tristate_controller_0_tcm_chipselect_n_out -> tristate_conduit_bridge_0:tcs_generic_tristate_controller_0_tcm_chipselect_n_out
	wire          tristate_conduit_pin_sharer_0_tcm_generic_tristate_controller_0_tcm_data_out_outen;                                   // tristate_conduit_pin_sharer_0:generic_tristate_controller_0_tcm_data_outen -> tristate_conduit_bridge_0:tcs_generic_tristate_controller_0_tcm_data_outen
	wire   [21:0] tristate_conduit_pin_sharer_0_tcm_generic_tristate_controller_0_tcm_address_out_out;                                  // tristate_conduit_pin_sharer_0:generic_tristate_controller_0_tcm_address_out -> tristate_conduit_bridge_0:tcs_generic_tristate_controller_0_tcm_address_out
	wire          generic_tristate_controller_0_tcm_chipselect_n_out;                                                                   // generic_tristate_controller_0:tcm_chipselect_n_out -> tristate_conduit_pin_sharer_0:tcs0_chipselect_n_out
	wire          generic_tristate_controller_0_tcm_grant;                                                                              // tristate_conduit_pin_sharer_0:tcs0_grant -> generic_tristate_controller_0:tcm_grant
	wire          generic_tristate_controller_0_tcm_data_outen;                                                                         // generic_tristate_controller_0:tcm_data_outen -> tristate_conduit_pin_sharer_0:tcs0_data_outen
	wire          generic_tristate_controller_0_tcm_request;                                                                            // generic_tristate_controller_0:tcm_request -> tristate_conduit_pin_sharer_0:tcs0_request
	wire    [7:0] generic_tristate_controller_0_tcm_data_out;                                                                           // generic_tristate_controller_0:tcm_data_out -> tristate_conduit_pin_sharer_0:tcs0_data_out
	wire          generic_tristate_controller_0_tcm_write_n_out;                                                                        // generic_tristate_controller_0:tcm_write_n_out -> tristate_conduit_pin_sharer_0:tcs0_write_n_out
	wire   [21:0] generic_tristate_controller_0_tcm_address_out;                                                                        // generic_tristate_controller_0:tcm_address_out -> tristate_conduit_pin_sharer_0:tcs0_address_out
	wire    [7:0] generic_tristate_controller_0_tcm_data_in;                                                                            // tristate_conduit_pin_sharer_0:tcs0_data_in -> generic_tristate_controller_0:tcm_data_in
	wire          generic_tristate_controller_0_tcm_read_n_out;                                                                         // generic_tristate_controller_0:tcm_read_n_out -> tristate_conduit_pin_sharer_0:tcs0_read_n_out
	wire          nios2_qsys_0_instruction_master_waitrequest;                                                                          // nios2_qsys_0_instruction_master_translator:av_waitrequest -> nios2_qsys_0:i_waitrequest
	wire   [24:0] nios2_qsys_0_instruction_master_address;                                                                              // nios2_qsys_0:i_address -> nios2_qsys_0_instruction_master_translator:av_address
	wire          nios2_qsys_0_instruction_master_read;                                                                                 // nios2_qsys_0:i_read -> nios2_qsys_0_instruction_master_translator:av_read
	wire   [31:0] nios2_qsys_0_instruction_master_readdata;                                                                             // nios2_qsys_0_instruction_master_translator:av_readdata -> nios2_qsys_0:i_readdata
	wire          nios2_qsys_0_instruction_master_readdatavalid;                                                                        // nios2_qsys_0_instruction_master_translator:av_readdatavalid -> nios2_qsys_0:i_readdatavalid
	wire          nios2_qsys_0_data_master_waitrequest;                                                                                 // nios2_qsys_0_data_master_translator:av_waitrequest -> nios2_qsys_0:d_waitrequest
	wire   [31:0] nios2_qsys_0_data_master_writedata;                                                                                   // nios2_qsys_0:d_writedata -> nios2_qsys_0_data_master_translator:av_writedata
	wire   [24:0] nios2_qsys_0_data_master_address;                                                                                     // nios2_qsys_0:d_address -> nios2_qsys_0_data_master_translator:av_address
	wire          nios2_qsys_0_data_master_write;                                                                                       // nios2_qsys_0:d_write -> nios2_qsys_0_data_master_translator:av_write
	wire          nios2_qsys_0_data_master_read;                                                                                        // nios2_qsys_0:d_read -> nios2_qsys_0_data_master_translator:av_read
	wire   [31:0] nios2_qsys_0_data_master_readdata;                                                                                    // nios2_qsys_0_data_master_translator:av_readdata -> nios2_qsys_0:d_readdata
	wire          nios2_qsys_0_data_master_debugaccess;                                                                                 // nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> nios2_qsys_0_data_master_translator:av_debugaccess
	wire          nios2_qsys_0_data_master_readdatavalid;                                                                               // nios2_qsys_0_data_master_translator:av_readdatavalid -> nios2_qsys_0:d_readdatavalid
	wire    [3:0] nios2_qsys_0_data_master_byteenable;                                                                                  // nios2_qsys_0:d_byteenable -> nios2_qsys_0_data_master_translator:av_byteenable
	wire   [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                              // nios2_qsys_0_jtag_debug_module_translator:av_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	wire    [8:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_address;                                                // nios2_qsys_0_jtag_debug_module_translator:av_address -> nios2_qsys_0:jtag_debug_module_address
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                                             // nios2_qsys_0_jtag_debug_module_translator:av_chipselect -> nios2_qsys_0:jtag_debug_module_select
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_write;                                                  // nios2_qsys_0_jtag_debug_module_translator:av_write -> nios2_qsys_0:jtag_debug_module_write
	wire   [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                               // nios2_qsys_0:jtag_debug_module_readdata -> nios2_qsys_0_jtag_debug_module_translator:av_readdata
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                                          // nios2_qsys_0_jtag_debug_module_translator:av_begintransfer -> nios2_qsys_0:jtag_debug_module_begintransfer
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                            // nios2_qsys_0_jtag_debug_module_translator:av_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	wire    [3:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                             // nios2_qsys_0_jtag_debug_module_translator:av_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata;                                                         // onchip_memory2_0_s1_translator:av_writedata -> onchip_memory2_0:writedata
	wire   [11:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_address;                                                           // onchip_memory2_0_s1_translator:av_address -> onchip_memory2_0:address
	wire          onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect;                                                        // onchip_memory2_0_s1_translator:av_chipselect -> onchip_memory2_0:chipselect
	wire          onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken;                                                             // onchip_memory2_0_s1_translator:av_clken -> onchip_memory2_0:clken
	wire          onchip_memory2_0_s1_translator_avalon_anti_slave_0_write;                                                             // onchip_memory2_0_s1_translator:av_write -> onchip_memory2_0:write
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata;                                                          // onchip_memory2_0:readdata -> onchip_memory2_0_s1_translator:av_readdata
	wire    [3:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable;                                                        // onchip_memory2_0_s1_translator:av_byteenable -> onchip_memory2_0:byteenable
	wire          sdram_0_s1_translator_avalon_anti_slave_0_waitrequest;                                                                // sdram_0:za_waitrequest -> sdram_0_s1_translator:av_waitrequest
	wire   [15:0] sdram_0_s1_translator_avalon_anti_slave_0_writedata;                                                                  // sdram_0_s1_translator:av_writedata -> sdram_0:az_data
	wire   [21:0] sdram_0_s1_translator_avalon_anti_slave_0_address;                                                                    // sdram_0_s1_translator:av_address -> sdram_0:az_addr
	wire          sdram_0_s1_translator_avalon_anti_slave_0_chipselect;                                                                 // sdram_0_s1_translator:av_chipselect -> sdram_0:az_cs
	wire          sdram_0_s1_translator_avalon_anti_slave_0_write;                                                                      // sdram_0_s1_translator:av_write -> sdram_0:az_wr_n
	wire          sdram_0_s1_translator_avalon_anti_slave_0_read;                                                                       // sdram_0_s1_translator:av_read -> sdram_0:az_rd_n
	wire   [15:0] sdram_0_s1_translator_avalon_anti_slave_0_readdata;                                                                   // sdram_0:za_data -> sdram_0_s1_translator:av_readdata
	wire          sdram_0_s1_translator_avalon_anti_slave_0_readdatavalid;                                                              // sdram_0:za_valid -> sdram_0_s1_translator:av_readdatavalid
	wire    [1:0] sdram_0_s1_translator_avalon_anti_slave_0_byteenable;                                                                 // sdram_0_s1_translator:av_byteenable -> sdram_0:az_be_n
	wire   [15:0] sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_writedata;                                                    // sram_0_avalon_sram_slave_translator:av_writedata -> sram_0:writedata
	wire   [17:0] sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_address;                                                      // sram_0_avalon_sram_slave_translator:av_address -> sram_0:address
	wire          sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_write;                                                        // sram_0_avalon_sram_slave_translator:av_write -> sram_0:write
	wire          sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_read;                                                         // sram_0_avalon_sram_slave_translator:av_read -> sram_0:read
	wire   [15:0] sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_readdata;                                                     // sram_0:readdata -> sram_0_avalon_sram_slave_translator:av_readdata
	wire          sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid;                                                // sram_0:readdatavalid -> sram_0_avalon_sram_slave_translator:av_readdatavalid
	wire    [1:0] sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable;                                                   // sram_0_avalon_sram_slave_translator:av_byteenable -> sram_0:byteenable
	wire   [15:0] sd_card_spi_master_spi_control_port_translator_avalon_anti_slave_0_writedata;                                         // sd_card_spi_master_spi_control_port_translator:av_writedata -> sd_card_spi_master:data_from_cpu
	wire    [2:0] sd_card_spi_master_spi_control_port_translator_avalon_anti_slave_0_address;                                           // sd_card_spi_master_spi_control_port_translator:av_address -> sd_card_spi_master:mem_addr
	wire          sd_card_spi_master_spi_control_port_translator_avalon_anti_slave_0_chipselect;                                        // sd_card_spi_master_spi_control_port_translator:av_chipselect -> sd_card_spi_master:spi_select
	wire          sd_card_spi_master_spi_control_port_translator_avalon_anti_slave_0_write;                                             // sd_card_spi_master_spi_control_port_translator:av_write -> sd_card_spi_master:write_n
	wire          sd_card_spi_master_spi_control_port_translator_avalon_anti_slave_0_read;                                              // sd_card_spi_master_spi_control_port_translator:av_read -> sd_card_spi_master:read_n
	wire   [15:0] sd_card_spi_master_spi_control_port_translator_avalon_anti_slave_0_readdata;                                          // sd_card_spi_master:data_to_cpu -> sd_card_spi_master_spi_control_port_translator:av_readdata
	wire          generic_tristate_controller_0_uas_translator_avalon_anti_slave_0_waitrequest;                                         // generic_tristate_controller_0:uas_waitrequest -> generic_tristate_controller_0_uas_translator:av_waitrequest
	wire    [0:0] generic_tristate_controller_0_uas_translator_avalon_anti_slave_0_burstcount;                                          // generic_tristate_controller_0_uas_translator:av_burstcount -> generic_tristate_controller_0:uas_burstcount
	wire    [7:0] generic_tristate_controller_0_uas_translator_avalon_anti_slave_0_writedata;                                           // generic_tristate_controller_0_uas_translator:av_writedata -> generic_tristate_controller_0:uas_writedata
	wire   [21:0] generic_tristate_controller_0_uas_translator_avalon_anti_slave_0_address;                                             // generic_tristate_controller_0_uas_translator:av_address -> generic_tristate_controller_0:uas_address
	wire          generic_tristate_controller_0_uas_translator_avalon_anti_slave_0_lock;                                                // generic_tristate_controller_0_uas_translator:av_lock -> generic_tristate_controller_0:uas_lock
	wire          generic_tristate_controller_0_uas_translator_avalon_anti_slave_0_write;                                               // generic_tristate_controller_0_uas_translator:av_write -> generic_tristate_controller_0:uas_write
	wire          generic_tristate_controller_0_uas_translator_avalon_anti_slave_0_read;                                                // generic_tristate_controller_0_uas_translator:av_read -> generic_tristate_controller_0:uas_read
	wire    [7:0] generic_tristate_controller_0_uas_translator_avalon_anti_slave_0_readdata;                                            // generic_tristate_controller_0:uas_readdata -> generic_tristate_controller_0_uas_translator:av_readdata
	wire          generic_tristate_controller_0_uas_translator_avalon_anti_slave_0_debugaccess;                                         // generic_tristate_controller_0_uas_translator:av_debugaccess -> generic_tristate_controller_0:uas_debugaccess
	wire          generic_tristate_controller_0_uas_translator_avalon_anti_slave_0_readdatavalid;                                       // generic_tristate_controller_0:uas_readdatavalid -> generic_tristate_controller_0_uas_translator:av_readdatavalid
	wire    [0:0] generic_tristate_controller_0_uas_translator_avalon_anti_slave_0_byteenable;                                          // generic_tristate_controller_0_uas_translator:av_byteenable -> generic_tristate_controller_0:uas_byteenable
	wire   [31:0] altpll_0_pll_slave_translator_avalon_anti_slave_0_writedata;                                                          // altpll_0_pll_slave_translator:av_writedata -> altpll_0:writedata
	wire    [1:0] altpll_0_pll_slave_translator_avalon_anti_slave_0_address;                                                            // altpll_0_pll_slave_translator:av_address -> altpll_0:address
	wire          altpll_0_pll_slave_translator_avalon_anti_slave_0_write;                                                              // altpll_0_pll_slave_translator:av_write -> altpll_0:write
	wire          altpll_0_pll_slave_translator_avalon_anti_slave_0_read;                                                               // altpll_0_pll_slave_translator:av_read -> altpll_0:read
	wire   [31:0] altpll_0_pll_slave_translator_avalon_anti_slave_0_readdata;                                                           // altpll_0:readdata -> altpll_0_pll_slave_translator:av_readdata
	wire    [0:0] sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_address;                                                    // sysid_qsys_0_control_slave_translator:av_address -> sysid_qsys_0:address
	wire   [31:0] sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_readdata;                                                   // sysid_qsys_0:readdata -> sysid_qsys_0_control_slave_translator:av_readdata
	wire   [15:0] timer_0_s1_translator_avalon_anti_slave_0_writedata;                                                                  // timer_0_s1_translator:av_writedata -> timer_0:writedata
	wire    [2:0] timer_0_s1_translator_avalon_anti_slave_0_address;                                                                    // timer_0_s1_translator:av_address -> timer_0:address
	wire          timer_0_s1_translator_avalon_anti_slave_0_chipselect;                                                                 // timer_0_s1_translator:av_chipselect -> timer_0:chipselect
	wire          timer_0_s1_translator_avalon_anti_slave_0_write;                                                                      // timer_0_s1_translator:av_write -> timer_0:write_n
	wire   [15:0] timer_0_s1_translator_avalon_anti_slave_0_readdata;                                                                   // timer_0:readdata -> timer_0_s1_translator:av_readdata
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                                             // jtag_uart_0:av_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                                               // jtag_uart_0_avalon_jtag_slave_translator:av_writedata -> jtag_uart_0:av_writedata
	wire    [0:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                                 // jtag_uart_0_avalon_jtag_slave_translator:av_address -> jtag_uart_0:av_address
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                                              // jtag_uart_0_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_0:av_chipselect
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                                   // jtag_uart_0_avalon_jtag_slave_translator:av_write -> jtag_uart_0:av_write_n
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                                    // jtag_uart_0_avalon_jtag_slave_translator:av_read -> jtag_uart_0:av_read_n
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                                                // jtag_uart_0:av_readdata -> jtag_uart_0_avalon_jtag_slave_translator:av_readdata
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_waitrequest;                                          // character_lcd_0:waitrequest -> character_lcd_0_avalon_lcd_slave_translator:av_waitrequest
	wire    [7:0] character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_writedata;                                            // character_lcd_0_avalon_lcd_slave_translator:av_writedata -> character_lcd_0:writedata
	wire    [0:0] character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_address;                                              // character_lcd_0_avalon_lcd_slave_translator:av_address -> character_lcd_0:address
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_chipselect;                                           // character_lcd_0_avalon_lcd_slave_translator:av_chipselect -> character_lcd_0:chipselect
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_write;                                                // character_lcd_0_avalon_lcd_slave_translator:av_write -> character_lcd_0:write
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_read;                                                 // character_lcd_0_avalon_lcd_slave_translator:av_read -> character_lcd_0:read
	wire    [7:0] character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_readdata;                                             // character_lcd_0:readdata -> character_lcd_0_avalon_lcd_slave_translator:av_readdata
	wire   [31:0] green_leds_s1_translator_avalon_anti_slave_0_writedata;                                                               // green_leds_s1_translator:av_writedata -> green_leds:writedata
	wire    [1:0] green_leds_s1_translator_avalon_anti_slave_0_address;                                                                 // green_leds_s1_translator:av_address -> green_leds:address
	wire          green_leds_s1_translator_avalon_anti_slave_0_chipselect;                                                              // green_leds_s1_translator:av_chipselect -> green_leds:chipselect
	wire          green_leds_s1_translator_avalon_anti_slave_0_write;                                                                   // green_leds_s1_translator:av_write -> green_leds:write_n
	wire   [31:0] green_leds_s1_translator_avalon_anti_slave_0_readdata;                                                                // green_leds:readdata -> green_leds_s1_translator:av_readdata
	wire    [1:0] switch_s1_translator_avalon_anti_slave_0_address;                                                                     // switch_s1_translator:av_address -> switch:address
	wire   [31:0] switch_s1_translator_avalon_anti_slave_0_readdata;                                                                    // switch:readdata -> switch_s1_translator:av_readdata
	wire   [31:0] audio_0_avalon_audio_slave_translator_avalon_anti_slave_0_writedata;                                                  // audio_0_avalon_audio_slave_translator:av_writedata -> audio_0:writedata
	wire    [1:0] audio_0_avalon_audio_slave_translator_avalon_anti_slave_0_address;                                                    // audio_0_avalon_audio_slave_translator:av_address -> audio_0:address
	wire          audio_0_avalon_audio_slave_translator_avalon_anti_slave_0_chipselect;                                                 // audio_0_avalon_audio_slave_translator:av_chipselect -> audio_0:chipselect
	wire          audio_0_avalon_audio_slave_translator_avalon_anti_slave_0_write;                                                      // audio_0_avalon_audio_slave_translator:av_write -> audio_0:write
	wire          audio_0_avalon_audio_slave_translator_avalon_anti_slave_0_read;                                                       // audio_0_avalon_audio_slave_translator:av_read -> audio_0:read
	wire   [31:0] audio_0_avalon_audio_slave_translator_avalon_anti_slave_0_readdata;                                                   // audio_0:readdata -> audio_0_avalon_audio_slave_translator:av_readdata
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_waitrequest;                           // audio_and_video_config_0:waitrequest -> audio_and_video_config_0_avalon_av_config_slave_translator:av_waitrequest
	wire   [31:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_writedata;                             // audio_and_video_config_0_avalon_av_config_slave_translator:av_writedata -> audio_and_video_config_0:writedata
	wire    [1:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_address;                               // audio_and_video_config_0_avalon_av_config_slave_translator:av_address -> audio_and_video_config_0:address
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_write;                                 // audio_and_video_config_0_avalon_av_config_slave_translator:av_write -> audio_and_video_config_0:write
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_read;                                  // audio_and_video_config_0_avalon_av_config_slave_translator:av_read -> audio_and_video_config_0:read
	wire   [31:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_readdata;                              // audio_and_video_config_0:readdata -> audio_and_video_config_0_avalon_av_config_slave_translator:av_readdata
	wire    [3:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_byteenable;                            // audio_and_video_config_0_avalon_av_config_slave_translator:av_byteenable -> audio_and_video_config_0:byteenable
	wire   [31:0] i2c_scl_s1_translator_avalon_anti_slave_0_writedata;                                                                  // I2C_SCL_s1_translator:av_writedata -> I2C_SCL:writedata
	wire    [1:0] i2c_scl_s1_translator_avalon_anti_slave_0_address;                                                                    // I2C_SCL_s1_translator:av_address -> I2C_SCL:address
	wire          i2c_scl_s1_translator_avalon_anti_slave_0_chipselect;                                                                 // I2C_SCL_s1_translator:av_chipselect -> I2C_SCL:chipselect
	wire          i2c_scl_s1_translator_avalon_anti_slave_0_write;                                                                      // I2C_SCL_s1_translator:av_write -> I2C_SCL:write_n
	wire   [31:0] i2c_scl_s1_translator_avalon_anti_slave_0_readdata;                                                                   // I2C_SCL:readdata -> I2C_SCL_s1_translator:av_readdata
	wire   [31:0] i2c_sda_s1_translator_avalon_anti_slave_0_writedata;                                                                  // I2C_SDA_s1_translator:av_writedata -> I2C_SDA:writedata
	wire    [1:0] i2c_sda_s1_translator_avalon_anti_slave_0_address;                                                                    // I2C_SDA_s1_translator:av_address -> I2C_SDA:address
	wire          i2c_sda_s1_translator_avalon_anti_slave_0_chipselect;                                                                 // I2C_SDA_s1_translator:av_chipselect -> I2C_SDA:chipselect
	wire          i2c_sda_s1_translator_avalon_anti_slave_0_write;                                                                      // I2C_SDA_s1_translator:av_write -> I2C_SDA:write_n
	wire   [31:0] i2c_sda_s1_translator_avalon_anti_slave_0_readdata;                                                                   // I2C_SDA:readdata -> I2C_SDA_s1_translator:av_readdata
	wire   [31:0] i2c_scl_2_s1_translator_avalon_anti_slave_0_writedata;                                                                // I2C_SCL_2_s1_translator:av_writedata -> I2C_SCL_2:writedata
	wire    [1:0] i2c_scl_2_s1_translator_avalon_anti_slave_0_address;                                                                  // I2C_SCL_2_s1_translator:av_address -> I2C_SCL_2:address
	wire          i2c_scl_2_s1_translator_avalon_anti_slave_0_chipselect;                                                               // I2C_SCL_2_s1_translator:av_chipselect -> I2C_SCL_2:chipselect
	wire          i2c_scl_2_s1_translator_avalon_anti_slave_0_write;                                                                    // I2C_SCL_2_s1_translator:av_write -> I2C_SCL_2:write_n
	wire   [31:0] i2c_scl_2_s1_translator_avalon_anti_slave_0_readdata;                                                                 // I2C_SCL_2:readdata -> I2C_SCL_2_s1_translator:av_readdata
	wire   [31:0] i2c_sda_2_s1_translator_avalon_anti_slave_0_writedata;                                                                // I2C_SDA_2_s1_translator:av_writedata -> I2C_SDA_2:writedata
	wire    [1:0] i2c_sda_2_s1_translator_avalon_anti_slave_0_address;                                                                  // I2C_SDA_2_s1_translator:av_address -> I2C_SDA_2:address
	wire          i2c_sda_2_s1_translator_avalon_anti_slave_0_chipselect;                                                               // I2C_SDA_2_s1_translator:av_chipselect -> I2C_SDA_2:chipselect
	wire          i2c_sda_2_s1_translator_avalon_anti_slave_0_write;                                                                    // I2C_SDA_2_s1_translator:av_write -> I2C_SDA_2:write_n
	wire   [31:0] i2c_sda_2_s1_translator_avalon_anti_slave_0_readdata;                                                                 // I2C_SDA_2:readdata -> I2C_SDA_2_s1_translator:av_readdata
	wire   [31:0] drum_out_s1_translator_avalon_anti_slave_0_writedata;                                                                 // drum_out_s1_translator:av_writedata -> drum_out:writedata
	wire    [1:0] drum_out_s1_translator_avalon_anti_slave_0_address;                                                                   // drum_out_s1_translator:av_address -> drum_out:address
	wire          drum_out_s1_translator_avalon_anti_slave_0_chipselect;                                                                // drum_out_s1_translator:av_chipselect -> drum_out:chipselect
	wire          drum_out_s1_translator_avalon_anti_slave_0_write;                                                                     // drum_out_s1_translator:av_write -> drum_out:write_n
	wire   [31:0] drum_out_s1_translator_avalon_anti_slave_0_readdata;                                                                  // drum_out:readdata -> drum_out_s1_translator:av_readdata
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_waitrequest;                                     // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_0_instruction_master_translator:uav_waitrequest
	wire    [2:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_burstcount;                                      // nios2_qsys_0_instruction_master_translator:uav_burstcount -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_writedata;                                       // nios2_qsys_0_instruction_master_translator:uav_writedata -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [24:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_address;                                         // nios2_qsys_0_instruction_master_translator:uav_address -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_lock;                                            // nios2_qsys_0_instruction_master_translator:uav_lock -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_write;                                           // nios2_qsys_0_instruction_master_translator:uav_write -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_read;                                            // nios2_qsys_0_instruction_master_translator:uav_read -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdata;                                        // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_0_instruction_master_translator:uav_readdata
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_debugaccess;                                     // nios2_qsys_0_instruction_master_translator:uav_debugaccess -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_byteenable;                                      // nios2_qsys_0_instruction_master_translator:uav_byteenable -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdatavalid;                                   // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_0_instruction_master_translator:uav_readdatavalid
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_waitrequest;                                            // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_0_data_master_translator:uav_waitrequest
	wire    [2:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_burstcount;                                             // nios2_qsys_0_data_master_translator:uav_burstcount -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_writedata;                                              // nios2_qsys_0_data_master_translator:uav_writedata -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [24:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_address;                                                // nios2_qsys_0_data_master_translator:uav_address -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_lock;                                                   // nios2_qsys_0_data_master_translator:uav_lock -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_write;                                                  // nios2_qsys_0_data_master_translator:uav_write -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_read;                                                   // nios2_qsys_0_data_master_translator:uav_read -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdata;                                               // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_0_data_master_translator:uav_readdata
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_debugaccess;                                            // nios2_qsys_0_data_master_translator:uav_debugaccess -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_byteenable;                                             // nios2_qsys_0_data_master_translator:uav_byteenable -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdatavalid;                                          // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_0_data_master_translator:uav_readdatavalid
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // nios2_qsys_0_jtag_debug_module_translator:uav_waitrequest -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> nios2_qsys_0_jtag_debug_module_translator:uav_burstcount
	wire   [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                                // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> nios2_qsys_0_jtag_debug_module_translator:uav_writedata
	wire   [24:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                                  // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> nios2_qsys_0_jtag_debug_module_translator:uav_address
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                                    // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> nios2_qsys_0_jtag_debug_module_translator:uav_write
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                                     // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> nios2_qsys_0_jtag_debug_module_translator:uav_lock
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                                     // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> nios2_qsys_0_jtag_debug_module_translator:uav_read
	wire   [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // nios2_qsys_0_jtag_debug_module_translator:uav_readdata -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // nios2_qsys_0_jtag_debug_module_translator:uav_readdatavalid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> nios2_qsys_0_jtag_debug_module_translator:uav_debugaccess
	wire    [3:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> nios2_qsys_0_jtag_debug_module_translator:uav_byteenable
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [102:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                              // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [102:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                         // onchip_memory2_0_s1_translator:uav_waitrequest -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                          // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> onchip_memory2_0_s1_translator:uav_burstcount
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                           // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> onchip_memory2_0_s1_translator:uav_writedata
	wire   [24:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                             // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> onchip_memory2_0_s1_translator:uav_address
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                               // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> onchip_memory2_0_s1_translator:uav_write
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> onchip_memory2_0_s1_translator:uav_lock
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> onchip_memory2_0_s1_translator:uav_read
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                            // onchip_memory2_0_s1_translator:uav_readdata -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                       // onchip_memory2_0_s1_translator:uav_readdatavalid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                         // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> onchip_memory2_0_s1_translator:uav_debugaccess
	wire    [3:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                          // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> onchip_memory2_0_s1_translator:uav_byteenable
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                  // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                        // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [102:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                         // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                        // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                               // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                     // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                             // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [102:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                      // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                     // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                   // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                    // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                   // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                  // sdram_0_s1_translator:uav_waitrequest -> sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [1:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                   // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sdram_0_s1_translator:uav_burstcount
	wire   [15:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                    // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sdram_0_s1_translator:uav_writedata
	wire   [24:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                      // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> sdram_0_s1_translator:uav_address
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                        // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> sdram_0_s1_translator:uav_write
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                         // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sdram_0_s1_translator:uav_lock
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                         // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> sdram_0_s1_translator:uav_read
	wire   [15:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                     // sdram_0_s1_translator:uav_readdata -> sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                // sdram_0_s1_translator:uav_readdatavalid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                  // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sdram_0_s1_translator:uav_debugaccess
	wire    [1:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                   // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sdram_0_s1_translator:uav_byteenable
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                           // sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                 // sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                         // sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [84:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                  // sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                 // sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                        // sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                              // sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                      // sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [84:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                               // sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                              // sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                            // sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [15:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                             // sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                            // sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // sram_0_avalon_sram_slave_translator:uav_waitrequest -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [1:0] sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sram_0_avalon_sram_slave_translator:uav_burstcount
	wire   [15:0] sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sram_0_avalon_sram_slave_translator:uav_writedata
	wire   [24:0] sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address;                                        // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_address -> sram_0_avalon_sram_slave_translator:uav_address
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write;                                          // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_write -> sram_0_avalon_sram_slave_translator:uav_write
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                           // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sram_0_avalon_sram_slave_translator:uav_lock
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read;                                           // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_read -> sram_0_avalon_sram_slave_translator:uav_read
	wire   [15:0] sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // sram_0_avalon_sram_slave_translator:uav_readdata -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // sram_0_avalon_sram_slave_translator:uav_readdatavalid -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sram_0_avalon_sram_slave_translator:uav_debugaccess
	wire    [1:0] sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sram_0_avalon_sram_slave_translator:uav_byteenable
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [84:0] sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [84:0] sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [15:0] sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest;                         // sd_card_spi_master_spi_control_port_translator:uav_waitrequest -> sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount;                          // sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:m0_burstcount -> sd_card_spi_master_spi_control_port_translator:uav_burstcount
	wire   [31:0] sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_m0_writedata;                           // sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:m0_writedata -> sd_card_spi_master_spi_control_port_translator:uav_writedata
	wire   [24:0] sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_m0_address;                             // sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:m0_address -> sd_card_spi_master_spi_control_port_translator:uav_address
	wire          sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_m0_write;                               // sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:m0_write -> sd_card_spi_master_spi_control_port_translator:uav_write
	wire          sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_m0_lock;                                // sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:m0_lock -> sd_card_spi_master_spi_control_port_translator:uav_lock
	wire          sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_m0_read;                                // sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:m0_read -> sd_card_spi_master_spi_control_port_translator:uav_read
	wire   [31:0] sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdata;                            // sd_card_spi_master_spi_control_port_translator:uav_readdata -> sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                       // sd_card_spi_master_spi_control_port_translator:uav_readdatavalid -> sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess;                         // sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sd_card_spi_master_spi_control_port_translator:uav_debugaccess
	wire    [3:0] sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable;                          // sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:m0_byteenable -> sd_card_spi_master_spi_control_port_translator:uav_byteenable
	wire          sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                  // sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid;                        // sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_valid -> sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                // sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [102:0] sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_data;                         // sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_data -> sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready;                        // sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;               // sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                     // sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;             // sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [102:0] sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                      // sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                     // sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                   // sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                    // sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                   // sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // generic_tristate_controller_0_uas_translator:uav_waitrequest -> generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire          generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:m0_burstcount -> generic_tristate_controller_0_uas_translator:uav_burstcount
	wire    [7:0] generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_m0_writedata;                             // generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:m0_writedata -> generic_tristate_controller_0_uas_translator:uav_writedata
	wire   [24:0] generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_m0_address;                               // generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:m0_address -> generic_tristate_controller_0_uas_translator:uav_address
	wire          generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_m0_write;                                 // generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:m0_write -> generic_tristate_controller_0_uas_translator:uav_write
	wire          generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_m0_lock;                                  // generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:m0_lock -> generic_tristate_controller_0_uas_translator:uav_lock
	wire          generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_m0_read;                                  // generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:m0_read -> generic_tristate_controller_0_uas_translator:uav_read
	wire    [7:0] generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_m0_readdata;                              // generic_tristate_controller_0_uas_translator:uav_readdata -> generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // generic_tristate_controller_0_uas_translator:uav_readdatavalid -> generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:m0_debugaccess -> generic_tristate_controller_0_uas_translator:uav_debugaccess
	wire          generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:m0_byteenable -> generic_tristate_controller_0_uas_translator:uav_byteenable
	wire          generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:rf_source_valid -> generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [75:0] generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rf_source_data;                           // generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:rf_source_data -> generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [75:0] generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:rf_sink_ready -> generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire    [7:0] generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                          // altpll_0_pll_slave_translator:uav_waitrequest -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                           // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> altpll_0_pll_slave_translator:uav_burstcount
	wire   [31:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                            // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> altpll_0_pll_slave_translator:uav_writedata
	wire   [24:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_address;                                              // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_address -> altpll_0_pll_slave_translator:uav_address
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_write;                                                // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_write -> altpll_0_pll_slave_translator:uav_write
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                                 // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_lock -> altpll_0_pll_slave_translator:uav_lock
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_read;                                                 // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_read -> altpll_0_pll_slave_translator:uav_read
	wire   [31:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                             // altpll_0_pll_slave_translator:uav_readdata -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                        // altpll_0_pll_slave_translator:uav_readdatavalid -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                          // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> altpll_0_pll_slave_translator:uav_debugaccess
	wire    [3:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                           // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> altpll_0_pll_slave_translator:uav_byteenable
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                   // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                                         // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                 // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [102:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                          // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                                         // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                      // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                              // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [102:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                       // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                      // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                    // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [31:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                     // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                    // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                                    // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                                     // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                                    // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // sysid_qsys_0_control_slave_translator:uav_waitrequest -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_qsys_0_control_slave_translator:uav_burstcount
	wire   [31:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_qsys_0_control_slave_translator:uav_writedata
	wire   [24:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                                      // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_qsys_0_control_slave_translator:uav_address
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                                        // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_qsys_0_control_slave_translator:uav_write
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                         // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_qsys_0_control_slave_translator:uav_lock
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                                         // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_qsys_0_control_slave_translator:uav_read
	wire   [31:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // sysid_qsys_0_control_slave_translator:uav_readdata -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // sysid_qsys_0_control_slave_translator:uav_readdatavalid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_qsys_0_control_slave_translator:uav_debugaccess
	wire    [3:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_qsys_0_control_slave_translator:uav_byteenable
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [102:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [102:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                  // timer_0_s1_translator:uav_waitrequest -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                   // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_0_s1_translator:uav_burstcount
	wire   [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                    // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_0_s1_translator:uav_writedata
	wire   [24:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                      // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_0_s1_translator:uav_address
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                        // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_0_s1_translator:uav_write
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                         // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_0_s1_translator:uav_lock
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                         // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_0_s1_translator:uav_read
	wire   [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                     // timer_0_s1_translator:uav_readdata -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                // timer_0_s1_translator:uav_readdatavalid -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                  // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_0_s1_translator:uav_debugaccess
	wire    [3:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                   // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_0_s1_translator:uav_byteenable
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                           // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                 // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                         // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [102:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                  // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                 // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                        // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                              // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                      // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [102:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                               // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                              // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                            // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                             // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                            // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // jtag_uart_0_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_0_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_0_avalon_jtag_slave_translator:uav_writedata
	wire   [24:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                                   // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_0_avalon_jtag_slave_translator:uav_address
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                                     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_0_avalon_jtag_slave_translator:uav_write
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                      // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_0_avalon_jtag_slave_translator:uav_lock
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                                      // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_0_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // jtag_uart_0_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // jtag_uart_0_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_0_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_0_avalon_jtag_slave_translator:uav_byteenable
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [102:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                               // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [102:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // character_lcd_0_avalon_lcd_slave_translator:uav_waitrequest -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> character_lcd_0_avalon_lcd_slave_translator:uav_burstcount
	wire    [7:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                              // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> character_lcd_0_avalon_lcd_slave_translator:uav_writedata
	wire   [24:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_address;                                // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_address -> character_lcd_0_avalon_lcd_slave_translator:uav_address
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_write;                                  // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_write -> character_lcd_0_avalon_lcd_slave_translator:uav_write
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                   // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_lock -> character_lcd_0_avalon_lcd_slave_translator:uav_lock
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_read;                                   // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_read -> character_lcd_0_avalon_lcd_slave_translator:uav_read
	wire    [7:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                               // character_lcd_0_avalon_lcd_slave_translator:uav_readdata -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // character_lcd_0_avalon_lcd_slave_translator:uav_readdatavalid -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> character_lcd_0_avalon_lcd_slave_translator:uav_debugaccess
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> character_lcd_0_avalon_lcd_slave_translator:uav_byteenable
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [75:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                            // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [75:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire    [7:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                               // green_leds_s1_translator:uav_waitrequest -> green_leds_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] green_leds_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                // green_leds_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> green_leds_s1_translator:uav_burstcount
	wire   [31:0] green_leds_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                 // green_leds_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> green_leds_s1_translator:uav_writedata
	wire   [24:0] green_leds_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                   // green_leds_s1_translator_avalon_universal_slave_0_agent:m0_address -> green_leds_s1_translator:uav_address
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                     // green_leds_s1_translator_avalon_universal_slave_0_agent:m0_write -> green_leds_s1_translator:uav_write
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                      // green_leds_s1_translator_avalon_universal_slave_0_agent:m0_lock -> green_leds_s1_translator:uav_lock
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                      // green_leds_s1_translator_avalon_universal_slave_0_agent:m0_read -> green_leds_s1_translator:uav_read
	wire   [31:0] green_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                  // green_leds_s1_translator:uav_readdata -> green_leds_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                             // green_leds_s1_translator:uav_readdatavalid -> green_leds_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                               // green_leds_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> green_leds_s1_translator:uav_debugaccess
	wire    [3:0] green_leds_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                // green_leds_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> green_leds_s1_translator:uav_byteenable
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                        // green_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                              // green_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                      // green_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [102:0] green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                               // green_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                              // green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> green_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                     // green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> green_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                           // green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> green_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                   // green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> green_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [102:0] green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                            // green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> green_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                           // green_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                         // green_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> green_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                          // green_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> green_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                         // green_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> green_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          switch_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                   // switch_s1_translator:uav_waitrequest -> switch_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] switch_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                    // switch_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> switch_s1_translator:uav_burstcount
	wire   [31:0] switch_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                     // switch_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> switch_s1_translator:uav_writedata
	wire   [24:0] switch_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                       // switch_s1_translator_avalon_universal_slave_0_agent:m0_address -> switch_s1_translator:uav_address
	wire          switch_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                         // switch_s1_translator_avalon_universal_slave_0_agent:m0_write -> switch_s1_translator:uav_write
	wire          switch_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                          // switch_s1_translator_avalon_universal_slave_0_agent:m0_lock -> switch_s1_translator:uav_lock
	wire          switch_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                          // switch_s1_translator_avalon_universal_slave_0_agent:m0_read -> switch_s1_translator:uav_read
	wire   [31:0] switch_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                      // switch_s1_translator:uav_readdata -> switch_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          switch_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                 // switch_s1_translator:uav_readdatavalid -> switch_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          switch_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                   // switch_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> switch_s1_translator:uav_debugaccess
	wire    [3:0] switch_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                    // switch_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> switch_s1_translator:uav_byteenable
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                            // switch_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                  // switch_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                          // switch_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [102:0] switch_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                   // switch_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                  // switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> switch_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                         // switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> switch_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                               // switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> switch_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                       // switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> switch_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [102:0] switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                                // switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> switch_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                               // switch_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                             // switch_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> switch_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                              // switch_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> switch_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                             // switch_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> switch_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // audio_0_avalon_audio_slave_translator:uav_waitrequest -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> audio_0_avalon_audio_slave_translator:uav_burstcount
	wire   [31:0] audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> audio_0_avalon_audio_slave_translator:uav_writedata
	wire   [24:0] audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_address;                                      // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_address -> audio_0_avalon_audio_slave_translator:uav_address
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_write;                                        // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_write -> audio_0_avalon_audio_slave_translator:uav_write
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                         // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_lock -> audio_0_avalon_audio_slave_translator:uav_lock
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_read;                                         // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_read -> audio_0_avalon_audio_slave_translator:uav_read
	wire   [31:0] audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // audio_0_avalon_audio_slave_translator:uav_readdata -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // audio_0_avalon_audio_slave_translator:uav_readdatavalid -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> audio_0_avalon_audio_slave_translator:uav_debugaccess
	wire    [3:0] audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> audio_0_avalon_audio_slave_translator:uav_byteenable
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [102:0] audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [102:0] audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [31:0] audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                            // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                             // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                            // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // audio_and_video_config_0_avalon_av_config_slave_translator:uav_waitrequest -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> audio_and_video_config_0_avalon_av_config_slave_translator:uav_burstcount
	wire   [31:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> audio_and_video_config_0_avalon_av_config_slave_translator:uav_writedata
	wire   [24:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_address -> audio_and_video_config_0_avalon_av_config_slave_translator:uav_address
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_write -> audio_and_video_config_0_avalon_av_config_slave_translator:uav_write
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_lock -> audio_and_video_config_0_avalon_av_config_slave_translator:uav_lock
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_read -> audio_and_video_config_0_avalon_av_config_slave_translator:uav_read
	wire   [31:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // audio_and_video_config_0_avalon_av_config_slave_translator:uav_readdata -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // audio_and_video_config_0_avalon_av_config_slave_translator:uav_readdatavalid -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> audio_and_video_config_0_avalon_av_config_slave_translator:uav_debugaccess
	wire    [3:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> audio_and_video_config_0_avalon_av_config_slave_translator:uav_byteenable
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [102:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [102:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [31:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;       // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;        // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;       // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                  // I2C_SCL_s1_translator:uav_waitrequest -> I2C_SCL_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                   // I2C_SCL_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> I2C_SCL_s1_translator:uav_burstcount
	wire   [31:0] i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                    // I2C_SCL_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> I2C_SCL_s1_translator:uav_writedata
	wire   [24:0] i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                      // I2C_SCL_s1_translator_avalon_universal_slave_0_agent:m0_address -> I2C_SCL_s1_translator:uav_address
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                        // I2C_SCL_s1_translator_avalon_universal_slave_0_agent:m0_write -> I2C_SCL_s1_translator:uav_write
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                         // I2C_SCL_s1_translator_avalon_universal_slave_0_agent:m0_lock -> I2C_SCL_s1_translator:uav_lock
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                         // I2C_SCL_s1_translator_avalon_universal_slave_0_agent:m0_read -> I2C_SCL_s1_translator:uav_read
	wire   [31:0] i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                     // I2C_SCL_s1_translator:uav_readdata -> I2C_SCL_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                // I2C_SCL_s1_translator:uav_readdatavalid -> I2C_SCL_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                  // I2C_SCL_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> I2C_SCL_s1_translator:uav_debugaccess
	wire    [3:0] i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                   // I2C_SCL_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> I2C_SCL_s1_translator:uav_byteenable
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                           // I2C_SCL_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> I2C_SCL_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                 // I2C_SCL_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> I2C_SCL_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                         // I2C_SCL_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> I2C_SCL_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [102:0] i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                  // I2C_SCL_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> I2C_SCL_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                 // I2C_SCL_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> I2C_SCL_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                        // I2C_SCL_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> I2C_SCL_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                              // I2C_SCL_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> I2C_SCL_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                      // I2C_SCL_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> I2C_SCL_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [102:0] i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                               // I2C_SCL_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> I2C_SCL_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                              // I2C_SCL_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> I2C_SCL_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                            // I2C_SCL_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> I2C_SCL_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                             // I2C_SCL_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> I2C_SCL_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                            // I2C_SCL_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> I2C_SCL_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                  // I2C_SDA_s1_translator:uav_waitrequest -> I2C_SDA_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                   // I2C_SDA_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> I2C_SDA_s1_translator:uav_burstcount
	wire   [31:0] i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                    // I2C_SDA_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> I2C_SDA_s1_translator:uav_writedata
	wire   [24:0] i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                      // I2C_SDA_s1_translator_avalon_universal_slave_0_agent:m0_address -> I2C_SDA_s1_translator:uav_address
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                        // I2C_SDA_s1_translator_avalon_universal_slave_0_agent:m0_write -> I2C_SDA_s1_translator:uav_write
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                         // I2C_SDA_s1_translator_avalon_universal_slave_0_agent:m0_lock -> I2C_SDA_s1_translator:uav_lock
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                         // I2C_SDA_s1_translator_avalon_universal_slave_0_agent:m0_read -> I2C_SDA_s1_translator:uav_read
	wire   [31:0] i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                     // I2C_SDA_s1_translator:uav_readdata -> I2C_SDA_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                // I2C_SDA_s1_translator:uav_readdatavalid -> I2C_SDA_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                  // I2C_SDA_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> I2C_SDA_s1_translator:uav_debugaccess
	wire    [3:0] i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                   // I2C_SDA_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> I2C_SDA_s1_translator:uav_byteenable
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                           // I2C_SDA_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> I2C_SDA_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                 // I2C_SDA_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> I2C_SDA_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                         // I2C_SDA_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> I2C_SDA_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [102:0] i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                  // I2C_SDA_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> I2C_SDA_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                 // I2C_SDA_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> I2C_SDA_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                        // I2C_SDA_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> I2C_SDA_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                              // I2C_SDA_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> I2C_SDA_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                      // I2C_SDA_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> I2C_SDA_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [102:0] i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                               // I2C_SDA_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> I2C_SDA_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                              // I2C_SDA_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> I2C_SDA_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                            // I2C_SDA_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> I2C_SDA_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                             // I2C_SDA_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> I2C_SDA_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                            // I2C_SDA_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> I2C_SDA_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                // I2C_SCL_2_s1_translator:uav_waitrequest -> I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                 // I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> I2C_SCL_2_s1_translator:uav_burstcount
	wire   [31:0] i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                  // I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> I2C_SCL_2_s1_translator:uav_writedata
	wire   [24:0] i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                    // I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:m0_address -> I2C_SCL_2_s1_translator:uav_address
	wire          i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                      // I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:m0_write -> I2C_SCL_2_s1_translator:uav_write
	wire          i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                       // I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:m0_lock -> I2C_SCL_2_s1_translator:uav_lock
	wire          i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                       // I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:m0_read -> I2C_SCL_2_s1_translator:uav_read
	wire   [31:0] i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                   // I2C_SCL_2_s1_translator:uav_readdata -> I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                              // I2C_SCL_2_s1_translator:uav_readdatavalid -> I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                // I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> I2C_SCL_2_s1_translator:uav_debugaccess
	wire    [3:0] i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                 // I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> I2C_SCL_2_s1_translator:uav_byteenable
	wire          i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                         // I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                               // I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                       // I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [102:0] i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                // I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                               // I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                      // I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                            // I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                    // I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [102:0] i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                             // I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                            // I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                          // I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                           // I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                          // I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                // I2C_SDA_2_s1_translator:uav_waitrequest -> I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                 // I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> I2C_SDA_2_s1_translator:uav_burstcount
	wire   [31:0] i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                  // I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> I2C_SDA_2_s1_translator:uav_writedata
	wire   [24:0] i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                    // I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:m0_address -> I2C_SDA_2_s1_translator:uav_address
	wire          i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                      // I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:m0_write -> I2C_SDA_2_s1_translator:uav_write
	wire          i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                       // I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:m0_lock -> I2C_SDA_2_s1_translator:uav_lock
	wire          i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                       // I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:m0_read -> I2C_SDA_2_s1_translator:uav_read
	wire   [31:0] i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                   // I2C_SDA_2_s1_translator:uav_readdata -> I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                              // I2C_SDA_2_s1_translator:uav_readdatavalid -> I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                // I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> I2C_SDA_2_s1_translator:uav_debugaccess
	wire    [3:0] i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                 // I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> I2C_SDA_2_s1_translator:uav_byteenable
	wire          i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                         // I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                               // I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                       // I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [102:0] i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                // I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                               // I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                      // I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                            // I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                    // I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [102:0] i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                             // I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                            // I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                          // I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                           // I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                          // I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          drum_out_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                 // drum_out_s1_translator:uav_waitrequest -> drum_out_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] drum_out_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                  // drum_out_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> drum_out_s1_translator:uav_burstcount
	wire   [31:0] drum_out_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                   // drum_out_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> drum_out_s1_translator:uav_writedata
	wire   [24:0] drum_out_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                     // drum_out_s1_translator_avalon_universal_slave_0_agent:m0_address -> drum_out_s1_translator:uav_address
	wire          drum_out_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                       // drum_out_s1_translator_avalon_universal_slave_0_agent:m0_write -> drum_out_s1_translator:uav_write
	wire          drum_out_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                        // drum_out_s1_translator_avalon_universal_slave_0_agent:m0_lock -> drum_out_s1_translator:uav_lock
	wire          drum_out_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                        // drum_out_s1_translator_avalon_universal_slave_0_agent:m0_read -> drum_out_s1_translator:uav_read
	wire   [31:0] drum_out_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                    // drum_out_s1_translator:uav_readdata -> drum_out_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          drum_out_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                               // drum_out_s1_translator:uav_readdatavalid -> drum_out_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          drum_out_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                 // drum_out_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> drum_out_s1_translator:uav_debugaccess
	wire    [3:0] drum_out_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                  // drum_out_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> drum_out_s1_translator:uav_byteenable
	wire          drum_out_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                          // drum_out_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> drum_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          drum_out_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                // drum_out_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> drum_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          drum_out_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                        // drum_out_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> drum_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [102:0] drum_out_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                 // drum_out_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> drum_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          drum_out_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                // drum_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> drum_out_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          drum_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                       // drum_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> drum_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          drum_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                             // drum_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> drum_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          drum_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                     // drum_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> drum_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [102:0] drum_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                              // drum_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> drum_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          drum_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                             // drum_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> drum_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          drum_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                           // drum_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> drum_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] drum_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                            // drum_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> drum_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          drum_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                           // drum_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> drum_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                            // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                                  // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                          // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [101:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                                   // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                                  // addr_router:sink_ready -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                                   // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_valid;                                         // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                                 // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [101:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_data;                                          // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_ready;                                         // addr_router_001:sink_ready -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                                    // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [101:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                                     // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router:sink_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                         // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                               // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                       // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [101:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                               // id_router_001:sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                  // sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                        // sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                // sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire   [83:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                         // sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                        // id_router_002:sink_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                          // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire   [83:0] sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data;                                           // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_003:sink_ready -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket;                         // sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire          sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rp_valid;                               // sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire          sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket;                       // sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [101:0] sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rp_data;                                // sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire          sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rp_ready;                               // id_router_004:sink_ready -> sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:rp_ready
	wire          generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire          generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rp_valid;                                 // generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire          generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire   [74:0] generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rp_data;                                  // generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire          generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_005:sink_ready -> generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:rp_ready
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                          // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                                // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                        // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [101:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_data;                                                 // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                                // id_router_006:sink_ready -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                        // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [101:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                                         // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_007:sink_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                  // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                        // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [101:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                         // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                        // id_router_008:sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire  [101:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                                      // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_009:sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                  // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire   [74:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_data;                                   // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_010:sink_ready -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                               // green_leds_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                     // green_leds_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                             // green_leds_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire  [101:0] green_leds_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                      // green_leds_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                     // id_router_011:sink_ready -> green_leds_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                   // switch_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                         // switch_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                 // switch_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	wire  [101:0] switch_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                          // switch_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                         // id_router_012:sink_ready -> switch_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                        // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	wire  [101:0] audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_data;                                         // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_013:sink_ready -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	wire  [101:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_014:sink_ready -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                  // I2C_SCL_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                        // I2C_SCL_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                // I2C_SCL_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	wire  [101:0] i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                         // I2C_SCL_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	wire          i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                        // id_router_015:sink_ready -> I2C_SCL_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                  // I2C_SDA_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_016:sink_endofpacket
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                        // I2C_SDA_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_016:sink_valid
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                // I2C_SDA_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_016:sink_startofpacket
	wire  [101:0] i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                         // I2C_SDA_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_016:sink_data
	wire          i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                        // id_router_016:sink_ready -> I2C_SDA_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                // I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_017:sink_endofpacket
	wire          i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                      // I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_017:sink_valid
	wire          i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                              // I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_017:sink_startofpacket
	wire  [101:0] i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                       // I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_017:sink_data
	wire          i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                      // id_router_017:sink_ready -> I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                // I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_018:sink_endofpacket
	wire          i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                      // I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_018:sink_valid
	wire          i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                              // I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_018:sink_startofpacket
	wire  [101:0] i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                       // I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_018:sink_data
	wire          i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                      // id_router_018:sink_ready -> I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          drum_out_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                 // drum_out_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_019:sink_endofpacket
	wire          drum_out_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                       // drum_out_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_019:sink_valid
	wire          drum_out_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                               // drum_out_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_019:sink_startofpacket
	wire  [101:0] drum_out_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                        // drum_out_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_019:sink_data
	wire          drum_out_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                       // id_router_019:sink_ready -> drum_out_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          addr_router_src_endofpacket;                                                                                          // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire          addr_router_src_valid;                                                                                                // addr_router:src_valid -> limiter:cmd_sink_valid
	wire          addr_router_src_startofpacket;                                                                                        // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [101:0] addr_router_src_data;                                                                                                 // addr_router:src_data -> limiter:cmd_sink_data
	wire   [19:0] addr_router_src_channel;                                                                                              // addr_router:src_channel -> limiter:cmd_sink_channel
	wire          addr_router_src_ready;                                                                                                // limiter:cmd_sink_ready -> addr_router:src_ready
	wire          limiter_rsp_src_endofpacket;                                                                                          // limiter:rsp_src_endofpacket -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_rsp_src_valid;                                                                                                // limiter:rsp_src_valid -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_rsp_src_startofpacket;                                                                                        // limiter:rsp_src_startofpacket -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [101:0] limiter_rsp_src_data;                                                                                                 // limiter:rsp_src_data -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [19:0] limiter_rsp_src_channel;                                                                                              // limiter:rsp_src_channel -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_rsp_src_ready;                                                                                                // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire          addr_router_001_src_endofpacket;                                                                                      // addr_router_001:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	wire          addr_router_001_src_valid;                                                                                            // addr_router_001:src_valid -> limiter_001:cmd_sink_valid
	wire          addr_router_001_src_startofpacket;                                                                                    // addr_router_001:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	wire  [101:0] addr_router_001_src_data;                                                                                             // addr_router_001:src_data -> limiter_001:cmd_sink_data
	wire   [19:0] addr_router_001_src_channel;                                                                                          // addr_router_001:src_channel -> limiter_001:cmd_sink_channel
	wire          addr_router_001_src_ready;                                                                                            // limiter_001:cmd_sink_ready -> addr_router_001:src_ready
	wire          limiter_001_rsp_src_endofpacket;                                                                                      // limiter_001:rsp_src_endofpacket -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_001_rsp_src_valid;                                                                                            // limiter_001:rsp_src_valid -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_001_rsp_src_startofpacket;                                                                                    // limiter_001:rsp_src_startofpacket -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [101:0] limiter_001_rsp_src_data;                                                                                             // limiter_001:rsp_src_data -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [19:0] limiter_001_rsp_src_channel;                                                                                          // limiter_001:rsp_src_channel -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_001_rsp_src_ready;                                                                                            // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_001:rsp_src_ready
	wire          burst_adapter_source0_endofpacket;                                                                                    // burst_adapter:source0_endofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_source0_valid;                                                                                          // burst_adapter:source0_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_source0_startofpacket;                                                                                  // burst_adapter:source0_startofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [83:0] burst_adapter_source0_data;                                                                                           // burst_adapter:source0_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_source0_ready;                                                                                          // sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire   [19:0] burst_adapter_source0_channel;                                                                                        // burst_adapter:source0_channel -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_001_source0_endofpacket;                                                                                // burst_adapter_001:source0_endofpacket -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_001_source0_valid;                                                                                      // burst_adapter_001:source0_valid -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_001_source0_startofpacket;                                                                              // burst_adapter_001:source0_startofpacket -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [83:0] burst_adapter_001_source0_data;                                                                                       // burst_adapter_001:source0_data -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_001_source0_ready;                                                                                      // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_001:source0_ready
	wire   [19:0] burst_adapter_001_source0_channel;                                                                                    // burst_adapter_001:source0_channel -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_002_source0_endofpacket;                                                                                // burst_adapter_002:source0_endofpacket -> generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_002_source0_valid;                                                                                      // burst_adapter_002:source0_valid -> generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_002_source0_startofpacket;                                                                              // burst_adapter_002:source0_startofpacket -> generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [74:0] burst_adapter_002_source0_data;                                                                                       // burst_adapter_002:source0_data -> generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_002_source0_ready;                                                                                      // generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_002:source0_ready
	wire   [19:0] burst_adapter_002_source0_channel;                                                                                    // burst_adapter_002:source0_channel -> generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_003_source0_endofpacket;                                                                                // burst_adapter_003:source0_endofpacket -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_003_source0_valid;                                                                                      // burst_adapter_003:source0_valid -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_003_source0_startofpacket;                                                                              // burst_adapter_003:source0_startofpacket -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [74:0] burst_adapter_003_source0_data;                                                                                       // burst_adapter_003:source0_data -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_003_source0_ready;                                                                                      // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_003:source0_ready
	wire   [19:0] burst_adapter_003_source0_channel;                                                                                    // burst_adapter_003:source0_channel -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rst_controller_reset_out_reset;                                                                                       // rst_controller:reset_out -> [I2C_SCL:reset_n, I2C_SCL_2:reset_n, I2C_SCL_2_s1_translator:reset, I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:reset, I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, I2C_SCL_s1_translator:reset, I2C_SCL_s1_translator_avalon_universal_slave_0_agent:reset, I2C_SCL_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, I2C_SDA:reset_n, I2C_SDA_2:reset_n, I2C_SDA_2_s1_translator:reset, I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:reset, I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, I2C_SDA_s1_translator:reset, I2C_SDA_s1_translator_avalon_universal_slave_0_agent:reset, I2C_SDA_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router:reset, addr_router_001:reset, burst_adapter:reset, burst_adapter_001:reset, burst_adapter_002:reset, burst_adapter_003:reset, character_lcd_0:reset, character_lcd_0_avalon_lcd_slave_translator:reset, character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:reset, character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, cmd_xbar_mux_003:reset, cmd_xbar_mux_004:reset, cmd_xbar_mux_005:reset, crosser:in_reset, crosser_001:in_reset, crosser_002:in_reset, crosser_003:out_reset, crosser_004:out_reset, crosser_005:out_reset, drum_out:reset_n, drum_out_s1_translator:reset, drum_out_s1_translator_avalon_universal_slave_0_agent:reset, drum_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, generic_tristate_controller_0:reset_reset, generic_tristate_controller_0_uas_translator:reset, generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent:reset, generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, green_leds:reset_n, green_leds_s1_translator:reset, green_leds_s1_translator_avalon_universal_slave_0_agent:reset, green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, id_router_011:reset, id_router_012:reset, id_router_015:reset, id_router_016:reset, id_router_017:reset, id_router_018:reset, id_router_019:reset, irq_mapper:reset, jtag_uart_0:rst_n, jtag_uart_0_avalon_jtag_slave_translator:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter:reset, limiter_001:reset, nios2_qsys_0:reset_n, nios2_qsys_0_data_master_translator:reset, nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_0_instruction_master_translator:reset, nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_0_jtag_debug_module_translator:reset, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, onchip_memory2_0:reset, onchip_memory2_0_s1_translator:reset, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:reset, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_015:reset, rsp_xbar_demux_016:reset, rsp_xbar_demux_017:reset, rsp_xbar_demux_018:reset, rsp_xbar_demux_019:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, sd_card_spi_master:reset_n, sd_card_spi_master_spi_control_port_translator:reset, sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:reset, sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sdram_0:reset_n, sdram_0_s1_translator:reset, sdram_0_s1_translator_avalon_universal_slave_0_agent:reset, sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sram_0:reset, sram_0_avalon_sram_slave_translator:reset, sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:reset, sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, switch:reset_n, switch_s1_translator:reset, switch_s1_translator_avalon_universal_slave_0_agent:reset, switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sysid_qsys_0:reset_n, sysid_qsys_0_control_slave_translator:reset, sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer_0:reset_n, timer_0_s1_translator:reset, timer_0_s1_translator_avalon_universal_slave_0_agent:reset, timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, tristate_conduit_bridge_0:reset, tristate_conduit_pin_sharer_0:reset_reset, up_clocks_0:reset, up_clocks_1:reset, width_adapter:reset, width_adapter_001:reset, width_adapter_002:reset, width_adapter_003:reset, width_adapter_004:reset, width_adapter_005:reset, width_adapter_006:reset, width_adapter_007:reset]
	wire          nios2_qsys_0_jtag_debug_module_reset_reset;                                                                           // nios2_qsys_0:jtag_debug_module_resetrequest -> [rst_controller:reset_in0, rst_controller_001:reset_in1, rst_controller_002:reset_in0]
	wire          rst_controller_001_reset_out_reset;                                                                                   // rst_controller_001:reset_out -> [altpll_0:reset, altpll_0_pll_slave_translator:reset, altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:reset, altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, crosser:out_reset, crosser_003:in_reset, id_router_006:reset, rsp_xbar_demux_006:reset]
	wire          rst_controller_002_reset_out_reset;                                                                                   // rst_controller_002:reset_out -> [audio_0:reset, audio_0_avalon_audio_slave_translator:reset, audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:reset, audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, audio_and_video_config_0:reset, audio_and_video_config_0_avalon_av_config_slave_translator:reset, audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:reset, audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, crosser_001:out_reset, crosser_002:out_reset, crosser_004:in_reset, crosser_005:in_reset, id_router_013:reset, id_router_014:reset, rsp_xbar_demux_013:reset, rsp_xbar_demux_014:reset]
	wire          cmd_xbar_demux_src0_endofpacket;                                                                                      // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                                            // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                                                    // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [101:0] cmd_xbar_demux_src0_data;                                                                                             // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire   [19:0] cmd_xbar_demux_src0_channel;                                                                                          // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire          cmd_xbar_demux_src0_ready;                                                                                            // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire          cmd_xbar_demux_src1_endofpacket;                                                                                      // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                                                            // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                                                    // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [101:0] cmd_xbar_demux_src1_data;                                                                                             // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire   [19:0] cmd_xbar_demux_src1_channel;                                                                                          // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire          cmd_xbar_demux_src1_ready;                                                                                            // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire          cmd_xbar_demux_src2_endofpacket;                                                                                      // cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire          cmd_xbar_demux_src2_valid;                                                                                            // cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	wire          cmd_xbar_demux_src2_startofpacket;                                                                                    // cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire  [101:0] cmd_xbar_demux_src2_data;                                                                                             // cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	wire   [19:0] cmd_xbar_demux_src2_channel;                                                                                          // cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	wire          cmd_xbar_demux_src2_ready;                                                                                            // cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	wire          cmd_xbar_demux_src3_endofpacket;                                                                                      // cmd_xbar_demux:src3_endofpacket -> cmd_xbar_mux_003:sink0_endofpacket
	wire          cmd_xbar_demux_src3_valid;                                                                                            // cmd_xbar_demux:src3_valid -> cmd_xbar_mux_003:sink0_valid
	wire          cmd_xbar_demux_src3_startofpacket;                                                                                    // cmd_xbar_demux:src3_startofpacket -> cmd_xbar_mux_003:sink0_startofpacket
	wire  [101:0] cmd_xbar_demux_src3_data;                                                                                             // cmd_xbar_demux:src3_data -> cmd_xbar_mux_003:sink0_data
	wire   [19:0] cmd_xbar_demux_src3_channel;                                                                                          // cmd_xbar_demux:src3_channel -> cmd_xbar_mux_003:sink0_channel
	wire          cmd_xbar_demux_src3_ready;                                                                                            // cmd_xbar_mux_003:sink0_ready -> cmd_xbar_demux:src3_ready
	wire          cmd_xbar_demux_src4_endofpacket;                                                                                      // cmd_xbar_demux:src4_endofpacket -> cmd_xbar_mux_004:sink0_endofpacket
	wire          cmd_xbar_demux_src4_valid;                                                                                            // cmd_xbar_demux:src4_valid -> cmd_xbar_mux_004:sink0_valid
	wire          cmd_xbar_demux_src4_startofpacket;                                                                                    // cmd_xbar_demux:src4_startofpacket -> cmd_xbar_mux_004:sink0_startofpacket
	wire  [101:0] cmd_xbar_demux_src4_data;                                                                                             // cmd_xbar_demux:src4_data -> cmd_xbar_mux_004:sink0_data
	wire   [19:0] cmd_xbar_demux_src4_channel;                                                                                          // cmd_xbar_demux:src4_channel -> cmd_xbar_mux_004:sink0_channel
	wire          cmd_xbar_demux_src4_ready;                                                                                            // cmd_xbar_mux_004:sink0_ready -> cmd_xbar_demux:src4_ready
	wire          cmd_xbar_demux_src5_endofpacket;                                                                                      // cmd_xbar_demux:src5_endofpacket -> cmd_xbar_mux_005:sink0_endofpacket
	wire          cmd_xbar_demux_src5_valid;                                                                                            // cmd_xbar_demux:src5_valid -> cmd_xbar_mux_005:sink0_valid
	wire          cmd_xbar_demux_src5_startofpacket;                                                                                    // cmd_xbar_demux:src5_startofpacket -> cmd_xbar_mux_005:sink0_startofpacket
	wire  [101:0] cmd_xbar_demux_src5_data;                                                                                             // cmd_xbar_demux:src5_data -> cmd_xbar_mux_005:sink0_data
	wire   [19:0] cmd_xbar_demux_src5_channel;                                                                                          // cmd_xbar_demux:src5_channel -> cmd_xbar_mux_005:sink0_channel
	wire          cmd_xbar_demux_src5_ready;                                                                                            // cmd_xbar_mux_005:sink0_ready -> cmd_xbar_demux:src5_ready
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                                                  // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                                                        // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                                                // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [101:0] cmd_xbar_demux_001_src0_data;                                                                                         // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire   [19:0] cmd_xbar_demux_001_src0_channel;                                                                                      // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                                                        // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire          cmd_xbar_demux_001_src1_endofpacket;                                                                                  // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire          cmd_xbar_demux_001_src1_valid;                                                                                        // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire          cmd_xbar_demux_001_src1_startofpacket;                                                                                // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [101:0] cmd_xbar_demux_001_src1_data;                                                                                         // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire   [19:0] cmd_xbar_demux_001_src1_channel;                                                                                      // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire          cmd_xbar_demux_001_src1_ready;                                                                                        // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire          cmd_xbar_demux_001_src2_endofpacket;                                                                                  // cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire          cmd_xbar_demux_001_src2_valid;                                                                                        // cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_002:sink1_valid
	wire          cmd_xbar_demux_001_src2_startofpacket;                                                                                // cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire  [101:0] cmd_xbar_demux_001_src2_data;                                                                                         // cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_002:sink1_data
	wire   [19:0] cmd_xbar_demux_001_src2_channel;                                                                                      // cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_002:sink1_channel
	wire          cmd_xbar_demux_001_src2_ready;                                                                                        // cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src2_ready
	wire          cmd_xbar_demux_001_src3_endofpacket;                                                                                  // cmd_xbar_demux_001:src3_endofpacket -> cmd_xbar_mux_003:sink1_endofpacket
	wire          cmd_xbar_demux_001_src3_valid;                                                                                        // cmd_xbar_demux_001:src3_valid -> cmd_xbar_mux_003:sink1_valid
	wire          cmd_xbar_demux_001_src3_startofpacket;                                                                                // cmd_xbar_demux_001:src3_startofpacket -> cmd_xbar_mux_003:sink1_startofpacket
	wire  [101:0] cmd_xbar_demux_001_src3_data;                                                                                         // cmd_xbar_demux_001:src3_data -> cmd_xbar_mux_003:sink1_data
	wire   [19:0] cmd_xbar_demux_001_src3_channel;                                                                                      // cmd_xbar_demux_001:src3_channel -> cmd_xbar_mux_003:sink1_channel
	wire          cmd_xbar_demux_001_src3_ready;                                                                                        // cmd_xbar_mux_003:sink1_ready -> cmd_xbar_demux_001:src3_ready
	wire          cmd_xbar_demux_001_src4_endofpacket;                                                                                  // cmd_xbar_demux_001:src4_endofpacket -> cmd_xbar_mux_004:sink1_endofpacket
	wire          cmd_xbar_demux_001_src4_valid;                                                                                        // cmd_xbar_demux_001:src4_valid -> cmd_xbar_mux_004:sink1_valid
	wire          cmd_xbar_demux_001_src4_startofpacket;                                                                                // cmd_xbar_demux_001:src4_startofpacket -> cmd_xbar_mux_004:sink1_startofpacket
	wire  [101:0] cmd_xbar_demux_001_src4_data;                                                                                         // cmd_xbar_demux_001:src4_data -> cmd_xbar_mux_004:sink1_data
	wire   [19:0] cmd_xbar_demux_001_src4_channel;                                                                                      // cmd_xbar_demux_001:src4_channel -> cmd_xbar_mux_004:sink1_channel
	wire          cmd_xbar_demux_001_src4_ready;                                                                                        // cmd_xbar_mux_004:sink1_ready -> cmd_xbar_demux_001:src4_ready
	wire          cmd_xbar_demux_001_src5_endofpacket;                                                                                  // cmd_xbar_demux_001:src5_endofpacket -> cmd_xbar_mux_005:sink1_endofpacket
	wire          cmd_xbar_demux_001_src5_valid;                                                                                        // cmd_xbar_demux_001:src5_valid -> cmd_xbar_mux_005:sink1_valid
	wire          cmd_xbar_demux_001_src5_startofpacket;                                                                                // cmd_xbar_demux_001:src5_startofpacket -> cmd_xbar_mux_005:sink1_startofpacket
	wire  [101:0] cmd_xbar_demux_001_src5_data;                                                                                         // cmd_xbar_demux_001:src5_data -> cmd_xbar_mux_005:sink1_data
	wire   [19:0] cmd_xbar_demux_001_src5_channel;                                                                                      // cmd_xbar_demux_001:src5_channel -> cmd_xbar_mux_005:sink1_channel
	wire          cmd_xbar_demux_001_src5_ready;                                                                                        // cmd_xbar_mux_005:sink1_ready -> cmd_xbar_demux_001:src5_ready
	wire          cmd_xbar_demux_001_src7_endofpacket;                                                                                  // cmd_xbar_demux_001:src7_endofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src7_valid;                                                                                        // cmd_xbar_demux_001:src7_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src7_startofpacket;                                                                                // cmd_xbar_demux_001:src7_startofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [101:0] cmd_xbar_demux_001_src7_data;                                                                                         // cmd_xbar_demux_001:src7_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [19:0] cmd_xbar_demux_001_src7_channel;                                                                                      // cmd_xbar_demux_001:src7_channel -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src8_endofpacket;                                                                                  // cmd_xbar_demux_001:src8_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src8_valid;                                                                                        // cmd_xbar_demux_001:src8_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src8_startofpacket;                                                                                // cmd_xbar_demux_001:src8_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [101:0] cmd_xbar_demux_001_src8_data;                                                                                         // cmd_xbar_demux_001:src8_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [19:0] cmd_xbar_demux_001_src8_channel;                                                                                      // cmd_xbar_demux_001:src8_channel -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src9_endofpacket;                                                                                  // cmd_xbar_demux_001:src9_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src9_valid;                                                                                        // cmd_xbar_demux_001:src9_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src9_startofpacket;                                                                                // cmd_xbar_demux_001:src9_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [101:0] cmd_xbar_demux_001_src9_data;                                                                                         // cmd_xbar_demux_001:src9_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [19:0] cmd_xbar_demux_001_src9_channel;                                                                                      // cmd_xbar_demux_001:src9_channel -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src10_endofpacket;                                                                                 // cmd_xbar_demux_001:src10_endofpacket -> width_adapter_006:in_endofpacket
	wire          cmd_xbar_demux_001_src10_valid;                                                                                       // cmd_xbar_demux_001:src10_valid -> width_adapter_006:in_valid
	wire          cmd_xbar_demux_001_src10_startofpacket;                                                                               // cmd_xbar_demux_001:src10_startofpacket -> width_adapter_006:in_startofpacket
	wire  [101:0] cmd_xbar_demux_001_src10_data;                                                                                        // cmd_xbar_demux_001:src10_data -> width_adapter_006:in_data
	wire   [19:0] cmd_xbar_demux_001_src10_channel;                                                                                     // cmd_xbar_demux_001:src10_channel -> width_adapter_006:in_channel
	wire          cmd_xbar_demux_001_src11_endofpacket;                                                                                 // cmd_xbar_demux_001:src11_endofpacket -> green_leds_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src11_valid;                                                                                       // cmd_xbar_demux_001:src11_valid -> green_leds_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src11_startofpacket;                                                                               // cmd_xbar_demux_001:src11_startofpacket -> green_leds_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [101:0] cmd_xbar_demux_001_src11_data;                                                                                        // cmd_xbar_demux_001:src11_data -> green_leds_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [19:0] cmd_xbar_demux_001_src11_channel;                                                                                     // cmd_xbar_demux_001:src11_channel -> green_leds_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src12_endofpacket;                                                                                 // cmd_xbar_demux_001:src12_endofpacket -> switch_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src12_valid;                                                                                       // cmd_xbar_demux_001:src12_valid -> switch_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src12_startofpacket;                                                                               // cmd_xbar_demux_001:src12_startofpacket -> switch_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [101:0] cmd_xbar_demux_001_src12_data;                                                                                        // cmd_xbar_demux_001:src12_data -> switch_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [19:0] cmd_xbar_demux_001_src12_channel;                                                                                     // cmd_xbar_demux_001:src12_channel -> switch_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src15_endofpacket;                                                                                 // cmd_xbar_demux_001:src15_endofpacket -> I2C_SCL_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src15_valid;                                                                                       // cmd_xbar_demux_001:src15_valid -> I2C_SCL_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src15_startofpacket;                                                                               // cmd_xbar_demux_001:src15_startofpacket -> I2C_SCL_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [101:0] cmd_xbar_demux_001_src15_data;                                                                                        // cmd_xbar_demux_001:src15_data -> I2C_SCL_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [19:0] cmd_xbar_demux_001_src15_channel;                                                                                     // cmd_xbar_demux_001:src15_channel -> I2C_SCL_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src16_endofpacket;                                                                                 // cmd_xbar_demux_001:src16_endofpacket -> I2C_SDA_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src16_valid;                                                                                       // cmd_xbar_demux_001:src16_valid -> I2C_SDA_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src16_startofpacket;                                                                               // cmd_xbar_demux_001:src16_startofpacket -> I2C_SDA_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [101:0] cmd_xbar_demux_001_src16_data;                                                                                        // cmd_xbar_demux_001:src16_data -> I2C_SDA_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [19:0] cmd_xbar_demux_001_src16_channel;                                                                                     // cmd_xbar_demux_001:src16_channel -> I2C_SDA_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src17_endofpacket;                                                                                 // cmd_xbar_demux_001:src17_endofpacket -> I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src17_valid;                                                                                       // cmd_xbar_demux_001:src17_valid -> I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src17_startofpacket;                                                                               // cmd_xbar_demux_001:src17_startofpacket -> I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [101:0] cmd_xbar_demux_001_src17_data;                                                                                        // cmd_xbar_demux_001:src17_data -> I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [19:0] cmd_xbar_demux_001_src17_channel;                                                                                     // cmd_xbar_demux_001:src17_channel -> I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src18_endofpacket;                                                                                 // cmd_xbar_demux_001:src18_endofpacket -> I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src18_valid;                                                                                       // cmd_xbar_demux_001:src18_valid -> I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src18_startofpacket;                                                                               // cmd_xbar_demux_001:src18_startofpacket -> I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [101:0] cmd_xbar_demux_001_src18_data;                                                                                        // cmd_xbar_demux_001:src18_data -> I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [19:0] cmd_xbar_demux_001_src18_channel;                                                                                     // cmd_xbar_demux_001:src18_channel -> I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src19_endofpacket;                                                                                 // cmd_xbar_demux_001:src19_endofpacket -> drum_out_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src19_valid;                                                                                       // cmd_xbar_demux_001:src19_valid -> drum_out_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src19_startofpacket;                                                                               // cmd_xbar_demux_001:src19_startofpacket -> drum_out_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [101:0] cmd_xbar_demux_001_src19_data;                                                                                        // cmd_xbar_demux_001:src19_data -> drum_out_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [19:0] cmd_xbar_demux_001_src19_channel;                                                                                     // cmd_xbar_demux_001:src19_channel -> drum_out_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rsp_xbar_demux_src0_endofpacket;                                                                                      // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                                            // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                                                    // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [101:0] rsp_xbar_demux_src0_data;                                                                                             // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [19:0] rsp_xbar_demux_src0_channel;                                                                                          // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire          rsp_xbar_demux_src0_ready;                                                                                            // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire          rsp_xbar_demux_src1_endofpacket;                                                                                      // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire          rsp_xbar_demux_src1_valid;                                                                                            // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire          rsp_xbar_demux_src1_startofpacket;                                                                                    // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [101:0] rsp_xbar_demux_src1_data;                                                                                             // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire   [19:0] rsp_xbar_demux_src1_channel;                                                                                          // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire          rsp_xbar_demux_src1_ready;                                                                                            // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                                                  // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                                                        // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                                                // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [101:0] rsp_xbar_demux_001_src0_data;                                                                                         // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire   [19:0] rsp_xbar_demux_001_src0_channel;                                                                                      // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                                                        // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire          rsp_xbar_demux_001_src1_endofpacket;                                                                                  // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire          rsp_xbar_demux_001_src1_valid;                                                                                        // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire          rsp_xbar_demux_001_src1_startofpacket;                                                                                // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [101:0] rsp_xbar_demux_001_src1_data;                                                                                         // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire   [19:0] rsp_xbar_demux_001_src1_channel;                                                                                      // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire          rsp_xbar_demux_001_src1_ready;                                                                                        // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                                                  // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                                                        // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                                                // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [101:0] rsp_xbar_demux_002_src0_data;                                                                                         // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire   [19:0] rsp_xbar_demux_002_src0_channel;                                                                                      // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                                                        // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire          rsp_xbar_demux_002_src1_endofpacket;                                                                                  // rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire          rsp_xbar_demux_002_src1_valid;                                                                                        // rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink2_valid
	wire          rsp_xbar_demux_002_src1_startofpacket;                                                                                // rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [101:0] rsp_xbar_demux_002_src1_data;                                                                                         // rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink2_data
	wire   [19:0] rsp_xbar_demux_002_src1_channel;                                                                                      // rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink2_channel
	wire          rsp_xbar_demux_002_src1_ready;                                                                                        // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src1_ready
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                                                  // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                                                        // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                                                // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	wire  [101:0] rsp_xbar_demux_003_src0_data;                                                                                         // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	wire   [19:0] rsp_xbar_demux_003_src0_channel;                                                                                      // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                                                        // rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire          rsp_xbar_demux_003_src1_endofpacket;                                                                                  // rsp_xbar_demux_003:src1_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire          rsp_xbar_demux_003_src1_valid;                                                                                        // rsp_xbar_demux_003:src1_valid -> rsp_xbar_mux_001:sink3_valid
	wire          rsp_xbar_demux_003_src1_startofpacket;                                                                                // rsp_xbar_demux_003:src1_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [101:0] rsp_xbar_demux_003_src1_data;                                                                                         // rsp_xbar_demux_003:src1_data -> rsp_xbar_mux_001:sink3_data
	wire   [19:0] rsp_xbar_demux_003_src1_channel;                                                                                      // rsp_xbar_demux_003:src1_channel -> rsp_xbar_mux_001:sink3_channel
	wire          rsp_xbar_demux_003_src1_ready;                                                                                        // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src1_ready
	wire          rsp_xbar_demux_004_src0_endofpacket;                                                                                  // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux:sink4_endofpacket
	wire          rsp_xbar_demux_004_src0_valid;                                                                                        // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux:sink4_valid
	wire          rsp_xbar_demux_004_src0_startofpacket;                                                                                // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux:sink4_startofpacket
	wire  [101:0] rsp_xbar_demux_004_src0_data;                                                                                         // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux:sink4_data
	wire   [19:0] rsp_xbar_demux_004_src0_channel;                                                                                      // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux:sink4_channel
	wire          rsp_xbar_demux_004_src0_ready;                                                                                        // rsp_xbar_mux:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire          rsp_xbar_demux_004_src1_endofpacket;                                                                                  // rsp_xbar_demux_004:src1_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire          rsp_xbar_demux_004_src1_valid;                                                                                        // rsp_xbar_demux_004:src1_valid -> rsp_xbar_mux_001:sink4_valid
	wire          rsp_xbar_demux_004_src1_startofpacket;                                                                                // rsp_xbar_demux_004:src1_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [101:0] rsp_xbar_demux_004_src1_data;                                                                                         // rsp_xbar_demux_004:src1_data -> rsp_xbar_mux_001:sink4_data
	wire   [19:0] rsp_xbar_demux_004_src1_channel;                                                                                      // rsp_xbar_demux_004:src1_channel -> rsp_xbar_mux_001:sink4_channel
	wire          rsp_xbar_demux_004_src1_ready;                                                                                        // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src1_ready
	wire          rsp_xbar_demux_005_src0_endofpacket;                                                                                  // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux:sink5_endofpacket
	wire          rsp_xbar_demux_005_src0_valid;                                                                                        // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux:sink5_valid
	wire          rsp_xbar_demux_005_src0_startofpacket;                                                                                // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux:sink5_startofpacket
	wire  [101:0] rsp_xbar_demux_005_src0_data;                                                                                         // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux:sink5_data
	wire   [19:0] rsp_xbar_demux_005_src0_channel;                                                                                      // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux:sink5_channel
	wire          rsp_xbar_demux_005_src0_ready;                                                                                        // rsp_xbar_mux:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire          rsp_xbar_demux_005_src1_endofpacket;                                                                                  // rsp_xbar_demux_005:src1_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire          rsp_xbar_demux_005_src1_valid;                                                                                        // rsp_xbar_demux_005:src1_valid -> rsp_xbar_mux_001:sink5_valid
	wire          rsp_xbar_demux_005_src1_startofpacket;                                                                                // rsp_xbar_demux_005:src1_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [101:0] rsp_xbar_demux_005_src1_data;                                                                                         // rsp_xbar_demux_005:src1_data -> rsp_xbar_mux_001:sink5_data
	wire   [19:0] rsp_xbar_demux_005_src1_channel;                                                                                      // rsp_xbar_demux_005:src1_channel -> rsp_xbar_mux_001:sink5_channel
	wire          rsp_xbar_demux_005_src1_ready;                                                                                        // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src1_ready
	wire          rsp_xbar_demux_007_src0_endofpacket;                                                                                  // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire          rsp_xbar_demux_007_src0_valid;                                                                                        // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink7_valid
	wire          rsp_xbar_demux_007_src0_startofpacket;                                                                                // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire  [101:0] rsp_xbar_demux_007_src0_data;                                                                                         // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink7_data
	wire   [19:0] rsp_xbar_demux_007_src0_channel;                                                                                      // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink7_channel
	wire          rsp_xbar_demux_007_src0_ready;                                                                                        // rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire          rsp_xbar_demux_008_src0_endofpacket;                                                                                  // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	wire          rsp_xbar_demux_008_src0_valid;                                                                                        // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_001:sink8_valid
	wire          rsp_xbar_demux_008_src0_startofpacket;                                                                                // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	wire  [101:0] rsp_xbar_demux_008_src0_data;                                                                                         // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_001:sink8_data
	wire   [19:0] rsp_xbar_demux_008_src0_channel;                                                                                      // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_001:sink8_channel
	wire          rsp_xbar_demux_008_src0_ready;                                                                                        // rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src0_ready
	wire          rsp_xbar_demux_009_src0_endofpacket;                                                                                  // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	wire          rsp_xbar_demux_009_src0_valid;                                                                                        // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_001:sink9_valid
	wire          rsp_xbar_demux_009_src0_startofpacket;                                                                                // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	wire  [101:0] rsp_xbar_demux_009_src0_data;                                                                                         // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_001:sink9_data
	wire   [19:0] rsp_xbar_demux_009_src0_channel;                                                                                      // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_001:sink9_channel
	wire          rsp_xbar_demux_009_src0_ready;                                                                                        // rsp_xbar_mux_001:sink9_ready -> rsp_xbar_demux_009:src0_ready
	wire          rsp_xbar_demux_010_src0_endofpacket;                                                                                  // rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux_001:sink10_endofpacket
	wire          rsp_xbar_demux_010_src0_valid;                                                                                        // rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux_001:sink10_valid
	wire          rsp_xbar_demux_010_src0_startofpacket;                                                                                // rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux_001:sink10_startofpacket
	wire  [101:0] rsp_xbar_demux_010_src0_data;                                                                                         // rsp_xbar_demux_010:src0_data -> rsp_xbar_mux_001:sink10_data
	wire   [19:0] rsp_xbar_demux_010_src0_channel;                                                                                      // rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux_001:sink10_channel
	wire          rsp_xbar_demux_010_src0_ready;                                                                                        // rsp_xbar_mux_001:sink10_ready -> rsp_xbar_demux_010:src0_ready
	wire          rsp_xbar_demux_011_src0_endofpacket;                                                                                  // rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux_001:sink11_endofpacket
	wire          rsp_xbar_demux_011_src0_valid;                                                                                        // rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux_001:sink11_valid
	wire          rsp_xbar_demux_011_src0_startofpacket;                                                                                // rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux_001:sink11_startofpacket
	wire  [101:0] rsp_xbar_demux_011_src0_data;                                                                                         // rsp_xbar_demux_011:src0_data -> rsp_xbar_mux_001:sink11_data
	wire   [19:0] rsp_xbar_demux_011_src0_channel;                                                                                      // rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux_001:sink11_channel
	wire          rsp_xbar_demux_011_src0_ready;                                                                                        // rsp_xbar_mux_001:sink11_ready -> rsp_xbar_demux_011:src0_ready
	wire          rsp_xbar_demux_012_src0_endofpacket;                                                                                  // rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux_001:sink12_endofpacket
	wire          rsp_xbar_demux_012_src0_valid;                                                                                        // rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux_001:sink12_valid
	wire          rsp_xbar_demux_012_src0_startofpacket;                                                                                // rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux_001:sink12_startofpacket
	wire  [101:0] rsp_xbar_demux_012_src0_data;                                                                                         // rsp_xbar_demux_012:src0_data -> rsp_xbar_mux_001:sink12_data
	wire   [19:0] rsp_xbar_demux_012_src0_channel;                                                                                      // rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux_001:sink12_channel
	wire          rsp_xbar_demux_012_src0_ready;                                                                                        // rsp_xbar_mux_001:sink12_ready -> rsp_xbar_demux_012:src0_ready
	wire          rsp_xbar_demux_015_src0_endofpacket;                                                                                  // rsp_xbar_demux_015:src0_endofpacket -> rsp_xbar_mux_001:sink15_endofpacket
	wire          rsp_xbar_demux_015_src0_valid;                                                                                        // rsp_xbar_demux_015:src0_valid -> rsp_xbar_mux_001:sink15_valid
	wire          rsp_xbar_demux_015_src0_startofpacket;                                                                                // rsp_xbar_demux_015:src0_startofpacket -> rsp_xbar_mux_001:sink15_startofpacket
	wire  [101:0] rsp_xbar_demux_015_src0_data;                                                                                         // rsp_xbar_demux_015:src0_data -> rsp_xbar_mux_001:sink15_data
	wire   [19:0] rsp_xbar_demux_015_src0_channel;                                                                                      // rsp_xbar_demux_015:src0_channel -> rsp_xbar_mux_001:sink15_channel
	wire          rsp_xbar_demux_015_src0_ready;                                                                                        // rsp_xbar_mux_001:sink15_ready -> rsp_xbar_demux_015:src0_ready
	wire          rsp_xbar_demux_016_src0_endofpacket;                                                                                  // rsp_xbar_demux_016:src0_endofpacket -> rsp_xbar_mux_001:sink16_endofpacket
	wire          rsp_xbar_demux_016_src0_valid;                                                                                        // rsp_xbar_demux_016:src0_valid -> rsp_xbar_mux_001:sink16_valid
	wire          rsp_xbar_demux_016_src0_startofpacket;                                                                                // rsp_xbar_demux_016:src0_startofpacket -> rsp_xbar_mux_001:sink16_startofpacket
	wire  [101:0] rsp_xbar_demux_016_src0_data;                                                                                         // rsp_xbar_demux_016:src0_data -> rsp_xbar_mux_001:sink16_data
	wire   [19:0] rsp_xbar_demux_016_src0_channel;                                                                                      // rsp_xbar_demux_016:src0_channel -> rsp_xbar_mux_001:sink16_channel
	wire          rsp_xbar_demux_016_src0_ready;                                                                                        // rsp_xbar_mux_001:sink16_ready -> rsp_xbar_demux_016:src0_ready
	wire          rsp_xbar_demux_017_src0_endofpacket;                                                                                  // rsp_xbar_demux_017:src0_endofpacket -> rsp_xbar_mux_001:sink17_endofpacket
	wire          rsp_xbar_demux_017_src0_valid;                                                                                        // rsp_xbar_demux_017:src0_valid -> rsp_xbar_mux_001:sink17_valid
	wire          rsp_xbar_demux_017_src0_startofpacket;                                                                                // rsp_xbar_demux_017:src0_startofpacket -> rsp_xbar_mux_001:sink17_startofpacket
	wire  [101:0] rsp_xbar_demux_017_src0_data;                                                                                         // rsp_xbar_demux_017:src0_data -> rsp_xbar_mux_001:sink17_data
	wire   [19:0] rsp_xbar_demux_017_src0_channel;                                                                                      // rsp_xbar_demux_017:src0_channel -> rsp_xbar_mux_001:sink17_channel
	wire          rsp_xbar_demux_017_src0_ready;                                                                                        // rsp_xbar_mux_001:sink17_ready -> rsp_xbar_demux_017:src0_ready
	wire          rsp_xbar_demux_018_src0_endofpacket;                                                                                  // rsp_xbar_demux_018:src0_endofpacket -> rsp_xbar_mux_001:sink18_endofpacket
	wire          rsp_xbar_demux_018_src0_valid;                                                                                        // rsp_xbar_demux_018:src0_valid -> rsp_xbar_mux_001:sink18_valid
	wire          rsp_xbar_demux_018_src0_startofpacket;                                                                                // rsp_xbar_demux_018:src0_startofpacket -> rsp_xbar_mux_001:sink18_startofpacket
	wire  [101:0] rsp_xbar_demux_018_src0_data;                                                                                         // rsp_xbar_demux_018:src0_data -> rsp_xbar_mux_001:sink18_data
	wire   [19:0] rsp_xbar_demux_018_src0_channel;                                                                                      // rsp_xbar_demux_018:src0_channel -> rsp_xbar_mux_001:sink18_channel
	wire          rsp_xbar_demux_018_src0_ready;                                                                                        // rsp_xbar_mux_001:sink18_ready -> rsp_xbar_demux_018:src0_ready
	wire          rsp_xbar_demux_019_src0_endofpacket;                                                                                  // rsp_xbar_demux_019:src0_endofpacket -> rsp_xbar_mux_001:sink19_endofpacket
	wire          rsp_xbar_demux_019_src0_valid;                                                                                        // rsp_xbar_demux_019:src0_valid -> rsp_xbar_mux_001:sink19_valid
	wire          rsp_xbar_demux_019_src0_startofpacket;                                                                                // rsp_xbar_demux_019:src0_startofpacket -> rsp_xbar_mux_001:sink19_startofpacket
	wire  [101:0] rsp_xbar_demux_019_src0_data;                                                                                         // rsp_xbar_demux_019:src0_data -> rsp_xbar_mux_001:sink19_data
	wire   [19:0] rsp_xbar_demux_019_src0_channel;                                                                                      // rsp_xbar_demux_019:src0_channel -> rsp_xbar_mux_001:sink19_channel
	wire          rsp_xbar_demux_019_src0_ready;                                                                                        // rsp_xbar_mux_001:sink19_ready -> rsp_xbar_demux_019:src0_ready
	wire          limiter_cmd_src_endofpacket;                                                                                          // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          limiter_cmd_src_startofpacket;                                                                                        // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [101:0] limiter_cmd_src_data;                                                                                                 // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire   [19:0] limiter_cmd_src_channel;                                                                                              // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire          limiter_cmd_src_ready;                                                                                                // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                                                         // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                                               // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                                                       // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [101:0] rsp_xbar_mux_src_data;                                                                                                // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire   [19:0] rsp_xbar_mux_src_channel;                                                                                             // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire          rsp_xbar_mux_src_ready;                                                                                               // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire          limiter_001_cmd_src_endofpacket;                                                                                      // limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          limiter_001_cmd_src_startofpacket;                                                                                    // limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [101:0] limiter_001_cmd_src_data;                                                                                             // limiter_001:cmd_src_data -> cmd_xbar_demux_001:sink_data
	wire   [19:0] limiter_001_cmd_src_channel;                                                                                          // limiter_001:cmd_src_channel -> cmd_xbar_demux_001:sink_channel
	wire          limiter_001_cmd_src_ready;                                                                                            // cmd_xbar_demux_001:sink_ready -> limiter_001:cmd_src_ready
	wire          rsp_xbar_mux_001_src_endofpacket;                                                                                     // rsp_xbar_mux_001:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	wire          rsp_xbar_mux_001_src_valid;                                                                                           // rsp_xbar_mux_001:src_valid -> limiter_001:rsp_sink_valid
	wire          rsp_xbar_mux_001_src_startofpacket;                                                                                   // rsp_xbar_mux_001:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	wire  [101:0] rsp_xbar_mux_001_src_data;                                                                                            // rsp_xbar_mux_001:src_data -> limiter_001:rsp_sink_data
	wire   [19:0] rsp_xbar_mux_001_src_channel;                                                                                         // rsp_xbar_mux_001:src_channel -> limiter_001:rsp_sink_channel
	wire          rsp_xbar_mux_001_src_ready;                                                                                           // limiter_001:rsp_sink_ready -> rsp_xbar_mux_001:src_ready
	wire          cmd_xbar_mux_src_endofpacket;                                                                                         // cmd_xbar_mux:src_endofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_src_valid;                                                                                               // cmd_xbar_mux:src_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_src_startofpacket;                                                                                       // cmd_xbar_mux:src_startofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [101:0] cmd_xbar_mux_src_data;                                                                                                // cmd_xbar_mux:src_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire   [19:0] cmd_xbar_mux_src_channel;                                                                                             // cmd_xbar_mux:src_channel -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_src_ready;                                                                                               // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire          id_router_src_endofpacket;                                                                                            // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                                                                  // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                                                          // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [101:0] id_router_src_data;                                                                                                   // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [19:0] id_router_src_channel;                                                                                                // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                                                                  // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          cmd_xbar_mux_001_src_endofpacket;                                                                                     // cmd_xbar_mux_001:src_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_001_src_valid;                                                                                           // cmd_xbar_mux_001:src_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_001_src_startofpacket;                                                                                   // cmd_xbar_mux_001:src_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [101:0] cmd_xbar_mux_001_src_data;                                                                                            // cmd_xbar_mux_001:src_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [19:0] cmd_xbar_mux_001_src_channel;                                                                                         // cmd_xbar_mux_001:src_channel -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_001_src_ready;                                                                                           // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	wire          id_router_001_src_endofpacket;                                                                                        // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          id_router_001_src_valid;                                                                                              // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire          id_router_001_src_startofpacket;                                                                                      // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [101:0] id_router_001_src_data;                                                                                               // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire   [19:0] id_router_001_src_channel;                                                                                            // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire          id_router_001_src_ready;                                                                                              // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire          cmd_xbar_mux_004_src_endofpacket;                                                                                     // cmd_xbar_mux_004:src_endofpacket -> sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_004_src_valid;                                                                                           // cmd_xbar_mux_004:src_valid -> sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_004_src_startofpacket;                                                                                   // cmd_xbar_mux_004:src_startofpacket -> sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [101:0] cmd_xbar_mux_004_src_data;                                                                                            // cmd_xbar_mux_004:src_data -> sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:cp_data
	wire   [19:0] cmd_xbar_mux_004_src_channel;                                                                                         // cmd_xbar_mux_004:src_channel -> sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_004_src_ready;                                                                                           // sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_004:src_ready
	wire          id_router_004_src_endofpacket;                                                                                        // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire          id_router_004_src_valid;                                                                                              // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire          id_router_004_src_startofpacket;                                                                                      // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [101:0] id_router_004_src_data;                                                                                               // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire   [19:0] id_router_004_src_channel;                                                                                            // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire          id_router_004_src_ready;                                                                                              // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire          crosser_out_ready;                                                                                                    // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:cp_ready -> crosser:out_ready
	wire          id_router_006_src_endofpacket;                                                                                        // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire          id_router_006_src_valid;                                                                                              // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire          id_router_006_src_startofpacket;                                                                                      // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [101:0] id_router_006_src_data;                                                                                               // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire   [19:0] id_router_006_src_channel;                                                                                            // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire          id_router_006_src_ready;                                                                                              // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire          cmd_xbar_demux_001_src7_ready;                                                                                        // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src7_ready
	wire          id_router_007_src_endofpacket;                                                                                        // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire          id_router_007_src_valid;                                                                                              // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire          id_router_007_src_startofpacket;                                                                                      // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [101:0] id_router_007_src_data;                                                                                               // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire   [19:0] id_router_007_src_channel;                                                                                            // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire          id_router_007_src_ready;                                                                                              // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire          cmd_xbar_demux_001_src8_ready;                                                                                        // timer_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src8_ready
	wire          id_router_008_src_endofpacket;                                                                                        // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire          id_router_008_src_valid;                                                                                              // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire          id_router_008_src_startofpacket;                                                                                      // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [101:0] id_router_008_src_data;                                                                                               // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire   [19:0] id_router_008_src_channel;                                                                                            // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire          id_router_008_src_ready;                                                                                              // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire          cmd_xbar_demux_001_src9_ready;                                                                                        // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src9_ready
	wire          id_router_009_src_endofpacket;                                                                                        // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire          id_router_009_src_valid;                                                                                              // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire          id_router_009_src_startofpacket;                                                                                      // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire  [101:0] id_router_009_src_data;                                                                                               // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire   [19:0] id_router_009_src_channel;                                                                                            // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire          id_router_009_src_ready;                                                                                              // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire          cmd_xbar_demux_001_src11_ready;                                                                                       // green_leds_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src11_ready
	wire          id_router_011_src_endofpacket;                                                                                        // id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire          id_router_011_src_valid;                                                                                              // id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	wire          id_router_011_src_startofpacket;                                                                                      // id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire  [101:0] id_router_011_src_data;                                                                                               // id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	wire   [19:0] id_router_011_src_channel;                                                                                            // id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	wire          id_router_011_src_ready;                                                                                              // rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	wire          cmd_xbar_demux_001_src12_ready;                                                                                       // switch_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src12_ready
	wire          id_router_012_src_endofpacket;                                                                                        // id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire          id_router_012_src_valid;                                                                                              // id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	wire          id_router_012_src_startofpacket;                                                                                      // id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire  [101:0] id_router_012_src_data;                                                                                               // id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	wire   [19:0] id_router_012_src_channel;                                                                                            // id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	wire          id_router_012_src_ready;                                                                                              // rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	wire          crosser_001_out_ready;                                                                                                // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_001:out_ready
	wire          id_router_013_src_endofpacket;                                                                                        // id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	wire          id_router_013_src_valid;                                                                                              // id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	wire          id_router_013_src_startofpacket;                                                                                      // id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	wire  [101:0] id_router_013_src_data;                                                                                               // id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	wire   [19:0] id_router_013_src_channel;                                                                                            // id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	wire          id_router_013_src_ready;                                                                                              // rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	wire          crosser_002_out_ready;                                                                                                // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_002:out_ready
	wire          id_router_014_src_endofpacket;                                                                                        // id_router_014:src_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	wire          id_router_014_src_valid;                                                                                              // id_router_014:src_valid -> rsp_xbar_demux_014:sink_valid
	wire          id_router_014_src_startofpacket;                                                                                      // id_router_014:src_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	wire  [101:0] id_router_014_src_data;                                                                                               // id_router_014:src_data -> rsp_xbar_demux_014:sink_data
	wire   [19:0] id_router_014_src_channel;                                                                                            // id_router_014:src_channel -> rsp_xbar_demux_014:sink_channel
	wire          id_router_014_src_ready;                                                                                              // rsp_xbar_demux_014:sink_ready -> id_router_014:src_ready
	wire          cmd_xbar_demux_001_src15_ready;                                                                                       // I2C_SCL_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src15_ready
	wire          id_router_015_src_endofpacket;                                                                                        // id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	wire          id_router_015_src_valid;                                                                                              // id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	wire          id_router_015_src_startofpacket;                                                                                      // id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	wire  [101:0] id_router_015_src_data;                                                                                               // id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	wire   [19:0] id_router_015_src_channel;                                                                                            // id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	wire          id_router_015_src_ready;                                                                                              // rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	wire          cmd_xbar_demux_001_src16_ready;                                                                                       // I2C_SDA_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src16_ready
	wire          id_router_016_src_endofpacket;                                                                                        // id_router_016:src_endofpacket -> rsp_xbar_demux_016:sink_endofpacket
	wire          id_router_016_src_valid;                                                                                              // id_router_016:src_valid -> rsp_xbar_demux_016:sink_valid
	wire          id_router_016_src_startofpacket;                                                                                      // id_router_016:src_startofpacket -> rsp_xbar_demux_016:sink_startofpacket
	wire  [101:0] id_router_016_src_data;                                                                                               // id_router_016:src_data -> rsp_xbar_demux_016:sink_data
	wire   [19:0] id_router_016_src_channel;                                                                                            // id_router_016:src_channel -> rsp_xbar_demux_016:sink_channel
	wire          id_router_016_src_ready;                                                                                              // rsp_xbar_demux_016:sink_ready -> id_router_016:src_ready
	wire          cmd_xbar_demux_001_src17_ready;                                                                                       // I2C_SCL_2_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src17_ready
	wire          id_router_017_src_endofpacket;                                                                                        // id_router_017:src_endofpacket -> rsp_xbar_demux_017:sink_endofpacket
	wire          id_router_017_src_valid;                                                                                              // id_router_017:src_valid -> rsp_xbar_demux_017:sink_valid
	wire          id_router_017_src_startofpacket;                                                                                      // id_router_017:src_startofpacket -> rsp_xbar_demux_017:sink_startofpacket
	wire  [101:0] id_router_017_src_data;                                                                                               // id_router_017:src_data -> rsp_xbar_demux_017:sink_data
	wire   [19:0] id_router_017_src_channel;                                                                                            // id_router_017:src_channel -> rsp_xbar_demux_017:sink_channel
	wire          id_router_017_src_ready;                                                                                              // rsp_xbar_demux_017:sink_ready -> id_router_017:src_ready
	wire          cmd_xbar_demux_001_src18_ready;                                                                                       // I2C_SDA_2_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src18_ready
	wire          id_router_018_src_endofpacket;                                                                                        // id_router_018:src_endofpacket -> rsp_xbar_demux_018:sink_endofpacket
	wire          id_router_018_src_valid;                                                                                              // id_router_018:src_valid -> rsp_xbar_demux_018:sink_valid
	wire          id_router_018_src_startofpacket;                                                                                      // id_router_018:src_startofpacket -> rsp_xbar_demux_018:sink_startofpacket
	wire  [101:0] id_router_018_src_data;                                                                                               // id_router_018:src_data -> rsp_xbar_demux_018:sink_data
	wire   [19:0] id_router_018_src_channel;                                                                                            // id_router_018:src_channel -> rsp_xbar_demux_018:sink_channel
	wire          id_router_018_src_ready;                                                                                              // rsp_xbar_demux_018:sink_ready -> id_router_018:src_ready
	wire          cmd_xbar_demux_001_src19_ready;                                                                                       // drum_out_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src19_ready
	wire          id_router_019_src_endofpacket;                                                                                        // id_router_019:src_endofpacket -> rsp_xbar_demux_019:sink_endofpacket
	wire          id_router_019_src_valid;                                                                                              // id_router_019:src_valid -> rsp_xbar_demux_019:sink_valid
	wire          id_router_019_src_startofpacket;                                                                                      // id_router_019:src_startofpacket -> rsp_xbar_demux_019:sink_startofpacket
	wire  [101:0] id_router_019_src_data;                                                                                               // id_router_019:src_data -> rsp_xbar_demux_019:sink_data
	wire   [19:0] id_router_019_src_channel;                                                                                            // id_router_019:src_channel -> rsp_xbar_demux_019:sink_channel
	wire          id_router_019_src_ready;                                                                                              // rsp_xbar_demux_019:sink_ready -> id_router_019:src_ready
	wire          cmd_xbar_mux_002_src_endofpacket;                                                                                     // cmd_xbar_mux_002:src_endofpacket -> width_adapter:in_endofpacket
	wire          cmd_xbar_mux_002_src_valid;                                                                                           // cmd_xbar_mux_002:src_valid -> width_adapter:in_valid
	wire          cmd_xbar_mux_002_src_startofpacket;                                                                                   // cmd_xbar_mux_002:src_startofpacket -> width_adapter:in_startofpacket
	wire  [101:0] cmd_xbar_mux_002_src_data;                                                                                            // cmd_xbar_mux_002:src_data -> width_adapter:in_data
	wire   [19:0] cmd_xbar_mux_002_src_channel;                                                                                         // cmd_xbar_mux_002:src_channel -> width_adapter:in_channel
	wire          cmd_xbar_mux_002_src_ready;                                                                                           // width_adapter:in_ready -> cmd_xbar_mux_002:src_ready
	wire          width_adapter_src_endofpacket;                                                                                        // width_adapter:out_endofpacket -> burst_adapter:sink0_endofpacket
	wire          width_adapter_src_valid;                                                                                              // width_adapter:out_valid -> burst_adapter:sink0_valid
	wire          width_adapter_src_startofpacket;                                                                                      // width_adapter:out_startofpacket -> burst_adapter:sink0_startofpacket
	wire   [83:0] width_adapter_src_data;                                                                                               // width_adapter:out_data -> burst_adapter:sink0_data
	wire          width_adapter_src_ready;                                                                                              // burst_adapter:sink0_ready -> width_adapter:out_ready
	wire   [19:0] width_adapter_src_channel;                                                                                            // width_adapter:out_channel -> burst_adapter:sink0_channel
	wire          id_router_002_src_endofpacket;                                                                                        // id_router_002:src_endofpacket -> width_adapter_001:in_endofpacket
	wire          id_router_002_src_valid;                                                                                              // id_router_002:src_valid -> width_adapter_001:in_valid
	wire          id_router_002_src_startofpacket;                                                                                      // id_router_002:src_startofpacket -> width_adapter_001:in_startofpacket
	wire   [83:0] id_router_002_src_data;                                                                                               // id_router_002:src_data -> width_adapter_001:in_data
	wire   [19:0] id_router_002_src_channel;                                                                                            // id_router_002:src_channel -> width_adapter_001:in_channel
	wire          id_router_002_src_ready;                                                                                              // width_adapter_001:in_ready -> id_router_002:src_ready
	wire          width_adapter_001_src_endofpacket;                                                                                    // width_adapter_001:out_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          width_adapter_001_src_valid;                                                                                          // width_adapter_001:out_valid -> rsp_xbar_demux_002:sink_valid
	wire          width_adapter_001_src_startofpacket;                                                                                  // width_adapter_001:out_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [101:0] width_adapter_001_src_data;                                                                                           // width_adapter_001:out_data -> rsp_xbar_demux_002:sink_data
	wire          width_adapter_001_src_ready;                                                                                          // rsp_xbar_demux_002:sink_ready -> width_adapter_001:out_ready
	wire   [19:0] width_adapter_001_src_channel;                                                                                        // width_adapter_001:out_channel -> rsp_xbar_demux_002:sink_channel
	wire          cmd_xbar_mux_003_src_endofpacket;                                                                                     // cmd_xbar_mux_003:src_endofpacket -> width_adapter_002:in_endofpacket
	wire          cmd_xbar_mux_003_src_valid;                                                                                           // cmd_xbar_mux_003:src_valid -> width_adapter_002:in_valid
	wire          cmd_xbar_mux_003_src_startofpacket;                                                                                   // cmd_xbar_mux_003:src_startofpacket -> width_adapter_002:in_startofpacket
	wire  [101:0] cmd_xbar_mux_003_src_data;                                                                                            // cmd_xbar_mux_003:src_data -> width_adapter_002:in_data
	wire   [19:0] cmd_xbar_mux_003_src_channel;                                                                                         // cmd_xbar_mux_003:src_channel -> width_adapter_002:in_channel
	wire          cmd_xbar_mux_003_src_ready;                                                                                           // width_adapter_002:in_ready -> cmd_xbar_mux_003:src_ready
	wire          width_adapter_002_src_endofpacket;                                                                                    // width_adapter_002:out_endofpacket -> burst_adapter_001:sink0_endofpacket
	wire          width_adapter_002_src_valid;                                                                                          // width_adapter_002:out_valid -> burst_adapter_001:sink0_valid
	wire          width_adapter_002_src_startofpacket;                                                                                  // width_adapter_002:out_startofpacket -> burst_adapter_001:sink0_startofpacket
	wire   [83:0] width_adapter_002_src_data;                                                                                           // width_adapter_002:out_data -> burst_adapter_001:sink0_data
	wire          width_adapter_002_src_ready;                                                                                          // burst_adapter_001:sink0_ready -> width_adapter_002:out_ready
	wire   [19:0] width_adapter_002_src_channel;                                                                                        // width_adapter_002:out_channel -> burst_adapter_001:sink0_channel
	wire          id_router_003_src_endofpacket;                                                                                        // id_router_003:src_endofpacket -> width_adapter_003:in_endofpacket
	wire          id_router_003_src_valid;                                                                                              // id_router_003:src_valid -> width_adapter_003:in_valid
	wire          id_router_003_src_startofpacket;                                                                                      // id_router_003:src_startofpacket -> width_adapter_003:in_startofpacket
	wire   [83:0] id_router_003_src_data;                                                                                               // id_router_003:src_data -> width_adapter_003:in_data
	wire   [19:0] id_router_003_src_channel;                                                                                            // id_router_003:src_channel -> width_adapter_003:in_channel
	wire          id_router_003_src_ready;                                                                                              // width_adapter_003:in_ready -> id_router_003:src_ready
	wire          width_adapter_003_src_endofpacket;                                                                                    // width_adapter_003:out_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          width_adapter_003_src_valid;                                                                                          // width_adapter_003:out_valid -> rsp_xbar_demux_003:sink_valid
	wire          width_adapter_003_src_startofpacket;                                                                                  // width_adapter_003:out_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [101:0] width_adapter_003_src_data;                                                                                           // width_adapter_003:out_data -> rsp_xbar_demux_003:sink_data
	wire          width_adapter_003_src_ready;                                                                                          // rsp_xbar_demux_003:sink_ready -> width_adapter_003:out_ready
	wire   [19:0] width_adapter_003_src_channel;                                                                                        // width_adapter_003:out_channel -> rsp_xbar_demux_003:sink_channel
	wire          cmd_xbar_mux_005_src_endofpacket;                                                                                     // cmd_xbar_mux_005:src_endofpacket -> width_adapter_004:in_endofpacket
	wire          cmd_xbar_mux_005_src_valid;                                                                                           // cmd_xbar_mux_005:src_valid -> width_adapter_004:in_valid
	wire          cmd_xbar_mux_005_src_startofpacket;                                                                                   // cmd_xbar_mux_005:src_startofpacket -> width_adapter_004:in_startofpacket
	wire  [101:0] cmd_xbar_mux_005_src_data;                                                                                            // cmd_xbar_mux_005:src_data -> width_adapter_004:in_data
	wire   [19:0] cmd_xbar_mux_005_src_channel;                                                                                         // cmd_xbar_mux_005:src_channel -> width_adapter_004:in_channel
	wire          cmd_xbar_mux_005_src_ready;                                                                                           // width_adapter_004:in_ready -> cmd_xbar_mux_005:src_ready
	wire          width_adapter_004_src_endofpacket;                                                                                    // width_adapter_004:out_endofpacket -> burst_adapter_002:sink0_endofpacket
	wire          width_adapter_004_src_valid;                                                                                          // width_adapter_004:out_valid -> burst_adapter_002:sink0_valid
	wire          width_adapter_004_src_startofpacket;                                                                                  // width_adapter_004:out_startofpacket -> burst_adapter_002:sink0_startofpacket
	wire   [74:0] width_adapter_004_src_data;                                                                                           // width_adapter_004:out_data -> burst_adapter_002:sink0_data
	wire          width_adapter_004_src_ready;                                                                                          // burst_adapter_002:sink0_ready -> width_adapter_004:out_ready
	wire   [19:0] width_adapter_004_src_channel;                                                                                        // width_adapter_004:out_channel -> burst_adapter_002:sink0_channel
	wire          id_router_005_src_endofpacket;                                                                                        // id_router_005:src_endofpacket -> width_adapter_005:in_endofpacket
	wire          id_router_005_src_valid;                                                                                              // id_router_005:src_valid -> width_adapter_005:in_valid
	wire          id_router_005_src_startofpacket;                                                                                      // id_router_005:src_startofpacket -> width_adapter_005:in_startofpacket
	wire   [74:0] id_router_005_src_data;                                                                                               // id_router_005:src_data -> width_adapter_005:in_data
	wire   [19:0] id_router_005_src_channel;                                                                                            // id_router_005:src_channel -> width_adapter_005:in_channel
	wire          id_router_005_src_ready;                                                                                              // width_adapter_005:in_ready -> id_router_005:src_ready
	wire          width_adapter_005_src_endofpacket;                                                                                    // width_adapter_005:out_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire          width_adapter_005_src_valid;                                                                                          // width_adapter_005:out_valid -> rsp_xbar_demux_005:sink_valid
	wire          width_adapter_005_src_startofpacket;                                                                                  // width_adapter_005:out_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [101:0] width_adapter_005_src_data;                                                                                           // width_adapter_005:out_data -> rsp_xbar_demux_005:sink_data
	wire          width_adapter_005_src_ready;                                                                                          // rsp_xbar_demux_005:sink_ready -> width_adapter_005:out_ready
	wire   [19:0] width_adapter_005_src_channel;                                                                                        // width_adapter_005:out_channel -> rsp_xbar_demux_005:sink_channel
	wire          cmd_xbar_demux_001_src10_ready;                                                                                       // width_adapter_006:in_ready -> cmd_xbar_demux_001:src10_ready
	wire          width_adapter_006_src_endofpacket;                                                                                    // width_adapter_006:out_endofpacket -> burst_adapter_003:sink0_endofpacket
	wire          width_adapter_006_src_valid;                                                                                          // width_adapter_006:out_valid -> burst_adapter_003:sink0_valid
	wire          width_adapter_006_src_startofpacket;                                                                                  // width_adapter_006:out_startofpacket -> burst_adapter_003:sink0_startofpacket
	wire   [74:0] width_adapter_006_src_data;                                                                                           // width_adapter_006:out_data -> burst_adapter_003:sink0_data
	wire          width_adapter_006_src_ready;                                                                                          // burst_adapter_003:sink0_ready -> width_adapter_006:out_ready
	wire   [19:0] width_adapter_006_src_channel;                                                                                        // width_adapter_006:out_channel -> burst_adapter_003:sink0_channel
	wire          id_router_010_src_endofpacket;                                                                                        // id_router_010:src_endofpacket -> width_adapter_007:in_endofpacket
	wire          id_router_010_src_valid;                                                                                              // id_router_010:src_valid -> width_adapter_007:in_valid
	wire          id_router_010_src_startofpacket;                                                                                      // id_router_010:src_startofpacket -> width_adapter_007:in_startofpacket
	wire   [74:0] id_router_010_src_data;                                                                                               // id_router_010:src_data -> width_adapter_007:in_data
	wire   [19:0] id_router_010_src_channel;                                                                                            // id_router_010:src_channel -> width_adapter_007:in_channel
	wire          id_router_010_src_ready;                                                                                              // width_adapter_007:in_ready -> id_router_010:src_ready
	wire          width_adapter_007_src_endofpacket;                                                                                    // width_adapter_007:out_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire          width_adapter_007_src_valid;                                                                                          // width_adapter_007:out_valid -> rsp_xbar_demux_010:sink_valid
	wire          width_adapter_007_src_startofpacket;                                                                                  // width_adapter_007:out_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire  [101:0] width_adapter_007_src_data;                                                                                           // width_adapter_007:out_data -> rsp_xbar_demux_010:sink_data
	wire          width_adapter_007_src_ready;                                                                                          // rsp_xbar_demux_010:sink_ready -> width_adapter_007:out_ready
	wire   [19:0] width_adapter_007_src_channel;                                                                                        // width_adapter_007:out_channel -> rsp_xbar_demux_010:sink_channel
	wire          crosser_out_endofpacket;                                                                                              // crosser:out_endofpacket -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_out_valid;                                                                                                    // crosser:out_valid -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_out_startofpacket;                                                                                            // crosser:out_startofpacket -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [101:0] crosser_out_data;                                                                                                     // crosser:out_data -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [19:0] crosser_out_channel;                                                                                                  // crosser:out_channel -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src6_endofpacket;                                                                                  // cmd_xbar_demux_001:src6_endofpacket -> crosser:in_endofpacket
	wire          cmd_xbar_demux_001_src6_valid;                                                                                        // cmd_xbar_demux_001:src6_valid -> crosser:in_valid
	wire          cmd_xbar_demux_001_src6_startofpacket;                                                                                // cmd_xbar_demux_001:src6_startofpacket -> crosser:in_startofpacket
	wire  [101:0] cmd_xbar_demux_001_src6_data;                                                                                         // cmd_xbar_demux_001:src6_data -> crosser:in_data
	wire   [19:0] cmd_xbar_demux_001_src6_channel;                                                                                      // cmd_xbar_demux_001:src6_channel -> crosser:in_channel
	wire          cmd_xbar_demux_001_src6_ready;                                                                                        // crosser:in_ready -> cmd_xbar_demux_001:src6_ready
	wire          crosser_001_out_endofpacket;                                                                                          // crosser_001:out_endofpacket -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_001_out_valid;                                                                                                // crosser_001:out_valid -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_001_out_startofpacket;                                                                                        // crosser_001:out_startofpacket -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [101:0] crosser_001_out_data;                                                                                                 // crosser_001:out_data -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [19:0] crosser_001_out_channel;                                                                                              // crosser_001:out_channel -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src13_endofpacket;                                                                                 // cmd_xbar_demux_001:src13_endofpacket -> crosser_001:in_endofpacket
	wire          cmd_xbar_demux_001_src13_valid;                                                                                       // cmd_xbar_demux_001:src13_valid -> crosser_001:in_valid
	wire          cmd_xbar_demux_001_src13_startofpacket;                                                                               // cmd_xbar_demux_001:src13_startofpacket -> crosser_001:in_startofpacket
	wire  [101:0] cmd_xbar_demux_001_src13_data;                                                                                        // cmd_xbar_demux_001:src13_data -> crosser_001:in_data
	wire   [19:0] cmd_xbar_demux_001_src13_channel;                                                                                     // cmd_xbar_demux_001:src13_channel -> crosser_001:in_channel
	wire          cmd_xbar_demux_001_src13_ready;                                                                                       // crosser_001:in_ready -> cmd_xbar_demux_001:src13_ready
	wire          crosser_002_out_endofpacket;                                                                                          // crosser_002:out_endofpacket -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_002_out_valid;                                                                                                // crosser_002:out_valid -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_002_out_startofpacket;                                                                                        // crosser_002:out_startofpacket -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [101:0] crosser_002_out_data;                                                                                                 // crosser_002:out_data -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [19:0] crosser_002_out_channel;                                                                                              // crosser_002:out_channel -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src14_endofpacket;                                                                                 // cmd_xbar_demux_001:src14_endofpacket -> crosser_002:in_endofpacket
	wire          cmd_xbar_demux_001_src14_valid;                                                                                       // cmd_xbar_demux_001:src14_valid -> crosser_002:in_valid
	wire          cmd_xbar_demux_001_src14_startofpacket;                                                                               // cmd_xbar_demux_001:src14_startofpacket -> crosser_002:in_startofpacket
	wire  [101:0] cmd_xbar_demux_001_src14_data;                                                                                        // cmd_xbar_demux_001:src14_data -> crosser_002:in_data
	wire   [19:0] cmd_xbar_demux_001_src14_channel;                                                                                     // cmd_xbar_demux_001:src14_channel -> crosser_002:in_channel
	wire          cmd_xbar_demux_001_src14_ready;                                                                                       // crosser_002:in_ready -> cmd_xbar_demux_001:src14_ready
	wire          crosser_003_out_endofpacket;                                                                                          // crosser_003:out_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire          crosser_003_out_valid;                                                                                                // crosser_003:out_valid -> rsp_xbar_mux_001:sink6_valid
	wire          crosser_003_out_startofpacket;                                                                                        // crosser_003:out_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [101:0] crosser_003_out_data;                                                                                                 // crosser_003:out_data -> rsp_xbar_mux_001:sink6_data
	wire   [19:0] crosser_003_out_channel;                                                                                              // crosser_003:out_channel -> rsp_xbar_mux_001:sink6_channel
	wire          crosser_003_out_ready;                                                                                                // rsp_xbar_mux_001:sink6_ready -> crosser_003:out_ready
	wire          rsp_xbar_demux_006_src0_endofpacket;                                                                                  // rsp_xbar_demux_006:src0_endofpacket -> crosser_003:in_endofpacket
	wire          rsp_xbar_demux_006_src0_valid;                                                                                        // rsp_xbar_demux_006:src0_valid -> crosser_003:in_valid
	wire          rsp_xbar_demux_006_src0_startofpacket;                                                                                // rsp_xbar_demux_006:src0_startofpacket -> crosser_003:in_startofpacket
	wire  [101:0] rsp_xbar_demux_006_src0_data;                                                                                         // rsp_xbar_demux_006:src0_data -> crosser_003:in_data
	wire   [19:0] rsp_xbar_demux_006_src0_channel;                                                                                      // rsp_xbar_demux_006:src0_channel -> crosser_003:in_channel
	wire          rsp_xbar_demux_006_src0_ready;                                                                                        // crosser_003:in_ready -> rsp_xbar_demux_006:src0_ready
	wire          crosser_004_out_endofpacket;                                                                                          // crosser_004:out_endofpacket -> rsp_xbar_mux_001:sink13_endofpacket
	wire          crosser_004_out_valid;                                                                                                // crosser_004:out_valid -> rsp_xbar_mux_001:sink13_valid
	wire          crosser_004_out_startofpacket;                                                                                        // crosser_004:out_startofpacket -> rsp_xbar_mux_001:sink13_startofpacket
	wire  [101:0] crosser_004_out_data;                                                                                                 // crosser_004:out_data -> rsp_xbar_mux_001:sink13_data
	wire   [19:0] crosser_004_out_channel;                                                                                              // crosser_004:out_channel -> rsp_xbar_mux_001:sink13_channel
	wire          crosser_004_out_ready;                                                                                                // rsp_xbar_mux_001:sink13_ready -> crosser_004:out_ready
	wire          rsp_xbar_demux_013_src0_endofpacket;                                                                                  // rsp_xbar_demux_013:src0_endofpacket -> crosser_004:in_endofpacket
	wire          rsp_xbar_demux_013_src0_valid;                                                                                        // rsp_xbar_demux_013:src0_valid -> crosser_004:in_valid
	wire          rsp_xbar_demux_013_src0_startofpacket;                                                                                // rsp_xbar_demux_013:src0_startofpacket -> crosser_004:in_startofpacket
	wire  [101:0] rsp_xbar_demux_013_src0_data;                                                                                         // rsp_xbar_demux_013:src0_data -> crosser_004:in_data
	wire   [19:0] rsp_xbar_demux_013_src0_channel;                                                                                      // rsp_xbar_demux_013:src0_channel -> crosser_004:in_channel
	wire          rsp_xbar_demux_013_src0_ready;                                                                                        // crosser_004:in_ready -> rsp_xbar_demux_013:src0_ready
	wire          crosser_005_out_endofpacket;                                                                                          // crosser_005:out_endofpacket -> rsp_xbar_mux_001:sink14_endofpacket
	wire          crosser_005_out_valid;                                                                                                // crosser_005:out_valid -> rsp_xbar_mux_001:sink14_valid
	wire          crosser_005_out_startofpacket;                                                                                        // crosser_005:out_startofpacket -> rsp_xbar_mux_001:sink14_startofpacket
	wire  [101:0] crosser_005_out_data;                                                                                                 // crosser_005:out_data -> rsp_xbar_mux_001:sink14_data
	wire   [19:0] crosser_005_out_channel;                                                                                              // crosser_005:out_channel -> rsp_xbar_mux_001:sink14_channel
	wire          crosser_005_out_ready;                                                                                                // rsp_xbar_mux_001:sink14_ready -> crosser_005:out_ready
	wire          rsp_xbar_demux_014_src0_endofpacket;                                                                                  // rsp_xbar_demux_014:src0_endofpacket -> crosser_005:in_endofpacket
	wire          rsp_xbar_demux_014_src0_valid;                                                                                        // rsp_xbar_demux_014:src0_valid -> crosser_005:in_valid
	wire          rsp_xbar_demux_014_src0_startofpacket;                                                                                // rsp_xbar_demux_014:src0_startofpacket -> crosser_005:in_startofpacket
	wire  [101:0] rsp_xbar_demux_014_src0_data;                                                                                         // rsp_xbar_demux_014:src0_data -> crosser_005:in_data
	wire   [19:0] rsp_xbar_demux_014_src0_channel;                                                                                      // rsp_xbar_demux_014:src0_channel -> crosser_005:in_channel
	wire          rsp_xbar_demux_014_src0_ready;                                                                                        // crosser_005:in_ready -> rsp_xbar_demux_014:src0_ready
	wire   [19:0] limiter_cmd_valid_data;                                                                                               // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire   [19:0] limiter_001_cmd_valid_data;                                                                                           // limiter_001:cmd_src_valid -> cmd_xbar_demux_001:sink_valid
	wire          irq_mapper_receiver0_irq;                                                                                             // timer_0:irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver1_irq;                                                                                             // jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	wire          irq_mapper_receiver2_irq;                                                                                             // sd_card_spi_master:irq -> irq_mapper:receiver2_irq
	wire   [31:0] nios2_qsys_0_d_irq_irq;                                                                                               // irq_mapper:sender_irq -> nios2_qsys_0:d_irq

	niosII_system_nios2_qsys_0 nios2_qsys_0 (
		.clk                                   (altpll_0_c1_clk),                                                             //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                             //                   reset_n.reset_n
		.d_address                             (nios2_qsys_0_data_master_address),                                            //               data_master.address
		.d_byteenable                          (nios2_qsys_0_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (nios2_qsys_0_data_master_read),                                               //                          .read
		.d_readdata                            (nios2_qsys_0_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (nios2_qsys_0_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (nios2_qsys_0_data_master_write),                                              //                          .write
		.d_writedata                           (nios2_qsys_0_data_master_writedata),                                          //                          .writedata
		.d_readdatavalid                       (nios2_qsys_0_data_master_readdatavalid),                                      //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (nios2_qsys_0_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (nios2_qsys_0_instruction_master_read),                                        //                          .read
		.i_readdata                            (nios2_qsys_0_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (nios2_qsys_0_instruction_master_waitrequest),                                 //                          .waitrequest
		.i_readdatavalid                       (nios2_qsys_0_instruction_master_readdatavalid),                               //                          .readdatavalid
		.d_irq                                 (nios2_qsys_0_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_qsys_0_jtag_debug_module_reset_reset),                                  //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.no_ci_readra                          ()                                                                             // custom_instruction_master.readra
	);

	niosII_system_onchip_memory2_0 onchip_memory2_0 (
		.clk        (altpll_0_c1_clk),                                               //   clk1.clk
		.address    (onchip_memory2_0_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (onchip_memory2_0_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset)                                 // reset1.reset
	);

	niosII_system_sysid_qsys_0 sysid_qsys_0 (
		.clock    (altpll_0_c1_clk),                                                    //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                                    //         reset.reset_n
		.readdata (sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_readdata), // control_slave.readdata
		.address  (sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_address)   //              .address
	);

	niosII_system_timer_0 timer_0 (
		.clk        (altpll_0_c1_clk),                                      //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      // reset.reset_n
		.address    (timer_0_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_0_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_0_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_0_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_0_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)                              //   irq.irq
	);

	niosII_system_jtag_uart_0 jtag_uart_0 (
		.clk            (altpll_0_c1_clk),                                                          //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                          //             reset.reset_n
		.av_chipselect  (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                                  //               irq.irq
	);

	niosII_system_character_lcd_0 character_lcd_0 (
		.clk         (altpll_0_c1_clk),                                                             //        clock_reset.clk
		.reset       (rst_controller_reset_out_reset),                                              //  clock_reset_reset.reset
		.address     (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_address),     //   avalon_lcd_slave.address
		.chipselect  (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_chipselect),  //                   .chipselect
		.read        (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_read),        //                   .read
		.write       (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_write),       //                   .write
		.writedata   (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_writedata),   //                   .writedata
		.readdata    (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_readdata),    //                   .readdata
		.waitrequest (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_waitrequest), //                   .waitrequest
		.LCD_DATA    (character_lcd_0_external_interface_DATA),                                     // external_interface.export
		.LCD_ON      (character_lcd_0_external_interface_ON),                                       //                   .export
		.LCD_BLON    (character_lcd_0_external_interface_BLON),                                     //                   .export
		.LCD_EN      (character_lcd_0_external_interface_EN),                                       //                   .export
		.LCD_RS      (character_lcd_0_external_interface_RS),                                       //                   .export
		.LCD_RW      (character_lcd_0_external_interface_RW)                                        //                   .export
	);

	niosII_system_green_leds green_leds (
		.clk        (altpll_0_c1_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                         //               reset.reset_n
		.address    (green_leds_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~green_leds_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (green_leds_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (green_leds_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (green_leds_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (green_leds_external_connection_export)                    // external_connection.export
	);

	niosII_system_switch switch (
		.clk      (altpll_0_c1_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address  (switch_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (switch_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (switch_external_connection_export)                  // external_connection.export
	);

	niosII_system_altpll_0 altpll_0 (
		.clk       (clk_clk),                                                     //       inclk_interface.clk
		.reset     (rst_controller_001_reset_out_reset),                          // inclk_interface_reset.reset
		.read      (altpll_0_pll_slave_translator_avalon_anti_slave_0_read),      //             pll_slave.read
		.write     (altpll_0_pll_slave_translator_avalon_anti_slave_0_write),     //                      .write
		.address   (altpll_0_pll_slave_translator_avalon_anti_slave_0_address),   //                      .address
		.readdata  (altpll_0_pll_slave_translator_avalon_anti_slave_0_readdata),  //                      .readdata
		.writedata (altpll_0_pll_slave_translator_avalon_anti_slave_0_writedata), //                      .writedata
		.c0        (altpll_0_c0_clk),                                             //                    c0.clk
		.c1        (altpll_0_c1_clk),                                             //                    c1.clk
		.areset    (),                                                            //        areset_conduit.export
		.locked    (),                                                            //        locked_conduit.export
		.phasedone ()                                                             //     phasedone_conduit.export
	);

	niosII_system_sdram_0 sdram_0 (
		.clk            (altpll_0_c1_clk),                                         //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                         // reset.reset_n
		.az_addr        (sdram_0_s1_translator_avalon_anti_slave_0_address),       //    s1.address
		.az_be_n        (~sdram_0_s1_translator_avalon_anti_slave_0_byteenable),   //      .byteenable_n
		.az_cs          (sdram_0_s1_translator_avalon_anti_slave_0_chipselect),    //      .chipselect
		.az_data        (sdram_0_s1_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.az_rd_n        (~sdram_0_s1_translator_avalon_anti_slave_0_read),         //      .read_n
		.az_wr_n        (~sdram_0_s1_translator_avalon_anti_slave_0_write),        //      .write_n
		.za_data        (sdram_0_s1_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.za_valid       (sdram_0_s1_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.za_waitrequest (sdram_0_s1_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_0_wire_addr),                                       //  wire.export
		.zs_ba          (sdram_0_wire_ba),                                         //      .export
		.zs_cas_n       (sdram_0_wire_cas_n),                                      //      .export
		.zs_cke         (sdram_0_wire_cke),                                        //      .export
		.zs_cs_n        (sdram_0_wire_cs_n),                                       //      .export
		.zs_dq          (sdram_0_wire_dq),                                         //      .export
		.zs_dqm         (sdram_0_wire_dqm),                                        //      .export
		.zs_ras_n       (sdram_0_wire_ras_n),                                      //      .export
		.zs_we_n        (sdram_0_wire_we_n)                                        //      .export
	);

	niosII_system_sram_0 sram_0 (
		.clk           (altpll_0_c1_clk),                                                       //        clock_reset.clk
		.reset         (rst_controller_reset_out_reset),                                        //  clock_reset_reset.reset
		.SRAM_DQ       (sram_0_external_interface_DQ),                                          // external_interface.export
		.SRAM_ADDR     (sram_0_external_interface_ADDR),                                        //                   .export
		.SRAM_LB_N     (sram_0_external_interface_LB_N),                                        //                   .export
		.SRAM_UB_N     (sram_0_external_interface_UB_N),                                        //                   .export
		.SRAM_CE_N     (sram_0_external_interface_CE_N),                                        //                   .export
		.SRAM_OE_N     (sram_0_external_interface_OE_N),                                        //                   .export
		.SRAM_WE_N     (sram_0_external_interface_WE_N),                                        //                   .export
		.address       (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_address),       //  avalon_sram_slave.address
		.byteenable    (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable),    //                   .byteenable
		.read          (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_read),          //                   .read
		.write         (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_write),         //                   .write
		.writedata     (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_writedata),     //                   .writedata
		.readdata      (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_readdata),      //                   .readdata
		.readdatavalid (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid)  //                   .readdatavalid
	);

	niosII_system_audio_0 audio_0 (
		.clk         (up_clocks_1_audio_clk_clk),                                            //        clock_reset.clk
		.reset       (rst_controller_002_reset_out_reset),                                   //  clock_reset_reset.reset
		.address     (audio_0_avalon_audio_slave_translator_avalon_anti_slave_0_address),    // avalon_audio_slave.address
		.chipselect  (audio_0_avalon_audio_slave_translator_avalon_anti_slave_0_chipselect), //                   .chipselect
		.read        (audio_0_avalon_audio_slave_translator_avalon_anti_slave_0_read),       //                   .read
		.write       (audio_0_avalon_audio_slave_translator_avalon_anti_slave_0_write),      //                   .write
		.writedata   (audio_0_avalon_audio_slave_translator_avalon_anti_slave_0_writedata),  //                   .writedata
		.readdata    (audio_0_avalon_audio_slave_translator_avalon_anti_slave_0_readdata),   //                   .readdata
		.irq         (),                                                                     //          interrupt.irq
		.AUD_ADCDAT  (audio_0_external_interface_ADCDAT),                                    // external_interface.export
		.AUD_ADCLRCK (audio_0_external_interface_ADCLRCK),                                   //                   .export
		.AUD_BCLK    (audio_0_external_interface_BCLK),                                      //                   .export
		.AUD_DACDAT  (audio_0_external_interface_DACDAT),                                    //                   .export
		.AUD_DACLRCK (audio_0_external_interface_DACLRCK)                                    //                   .export
	);

	niosII_system_audio_and_video_config_0 audio_and_video_config_0 (
		.clk         (up_clocks_1_audio_clk_clk),                                                                  //            clock_reset.clk
		.reset       (rst_controller_002_reset_out_reset),                                                         //      clock_reset_reset.reset
		.address     (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_address),     // avalon_av_config_slave.address
		.byteenable  (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_byteenable),  //                       .byteenable
		.read        (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_read),        //                       .read
		.write       (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_write),       //                       .write
		.writedata   (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_writedata),   //                       .writedata
		.readdata    (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_readdata),    //                       .readdata
		.waitrequest (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_waitrequest), //                       .waitrequest
		.I2C_SDAT    (audio_and_video_config_0_external_interface_SDAT),                                           //     external_interface.export
		.I2C_SCLK    (audio_and_video_config_0_external_interface_SCLK)                                            //                       .export
	);

	niosII_system_up_clocks_0 up_clocks_0 (
		.CLOCK_50    (altpll_0_c1_clk),                //       clk_in_primary.clk
		.reset       (rst_controller_reset_out_reset), // clk_in_primary_reset.reset
		.sys_clk     (),                               //              sys_clk.clk
		.sys_reset_n (),                               //        sys_clk_reset.reset_n
		.CLOCK_27    (clk_1_clk),                      //     clk_in_secondary.clk
		.AUD_CLK     (up_clocks_0_audio_clk_clk)       //            audio_clk.clk
	);

	niosII_system_up_clocks_0 up_clocks_1 (
		.CLOCK_50    (altpll_0_c1_clk),                //       clk_in_primary.clk
		.reset       (rst_controller_reset_out_reset), // clk_in_primary_reset.reset
		.sys_clk     (),                               //              sys_clk.clk
		.sys_reset_n (),                               //        sys_clk_reset.reset_n
		.CLOCK_27    (clk_1_clk),                      //     clk_in_secondary.clk
		.AUD_CLK     (up_clocks_1_audio_clk_clk)       //            audio_clk.clk
	);

	niosII_system_sd_card_spi_master sd_card_spi_master (
		.clk           (altpll_0_c1_clk),                                                               //              clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                                               //            reset.reset_n
		.data_from_cpu (sd_card_spi_master_spi_control_port_translator_avalon_anti_slave_0_writedata),  // spi_control_port.writedata
		.data_to_cpu   (sd_card_spi_master_spi_control_port_translator_avalon_anti_slave_0_readdata),   //                 .readdata
		.mem_addr      (sd_card_spi_master_spi_control_port_translator_avalon_anti_slave_0_address),    //                 .address
		.read_n        (~sd_card_spi_master_spi_control_port_translator_avalon_anti_slave_0_read),      //                 .read_n
		.spi_select    (sd_card_spi_master_spi_control_port_translator_avalon_anti_slave_0_chipselect), //                 .chipselect
		.write_n       (~sd_card_spi_master_spi_control_port_translator_avalon_anti_slave_0_write),     //                 .write_n
		.irq           (irq_mapper_receiver2_irq),                                                      //              irq.irq
		.MISO          (spi_0_external_MISO),                                                           //         external.export
		.MOSI          (spi_0_external_MOSI),                                                           //                 .export
		.SCLK          (spi_0_external_SCLK),                                                           //                 .export
		.SS_n          (spi_0_external_SS_n)                                                            //                 .export
	);

	niosII_system_I2C_SCL i2c_scl (
		.clk        (altpll_0_c1_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address    (i2c_scl_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~i2c_scl_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (i2c_scl_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (i2c_scl_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (i2c_scl_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (i2c_scl_external_connection_export)                    // external_connection.export
	);

	niosII_system_I2C_SDA i2c_sda (
		.clk        (altpll_0_c1_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address    (i2c_sda_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~i2c_sda_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (i2c_sda_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (i2c_sda_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (i2c_sda_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.bidir_port (i2c_sda_external_connection_export)                    // external_connection.export
	);

	niosII_system_I2C_SCL i2c_scl_2 (
		.clk        (altpll_0_c1_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                        //               reset.reset_n
		.address    (i2c_scl_2_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~i2c_scl_2_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (i2c_scl_2_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (i2c_scl_2_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (i2c_scl_2_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (i2c_scl_2_external_connection_export)                    // external_connection.export
	);

	niosII_system_I2C_SDA i2c_sda_2 (
		.clk        (altpll_0_c1_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                        //               reset.reset_n
		.address    (i2c_sda_2_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~i2c_sda_2_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (i2c_sda_2_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (i2c_sda_2_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (i2c_sda_2_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.bidir_port (i2c_sda_2_external_connection_export)                    // external_connection.export
	);

	niosII_system_drum_out drum_out (
		.clk        (altpll_0_c1_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                       //               reset.reset_n
		.address    (drum_out_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~drum_out_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (drum_out_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (drum_out_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (drum_out_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (drum_out_external_connection_export)                    // external_connection.export
	);

	niosII_system_generic_tristate_controller_0 #(
		.TCM_ADDRESS_W                  (22),
		.TCM_DATA_W                     (8),
		.TCM_BYTEENABLE_W               (1),
		.TCM_READ_WAIT                  (160),
		.TCM_WRITE_WAIT                 (160),
		.TCM_SETUP_WAIT                 (40),
		.TCM_DATA_HOLD                  (40),
		.TCM_TURNAROUND_TIME            (2),
		.TCM_TIMING_UNITS               (0),
		.TCM_READLATENCY                (2),
		.TCM_SYMBOLS_PER_WORD           (1),
		.USE_READDATA                   (1),
		.USE_WRITEDATA                  (1),
		.USE_READ                       (1),
		.USE_WRITE                      (1),
		.USE_BYTEENABLE                 (0),
		.USE_CHIPSELECT                 (1),
		.USE_LOCK                       (0),
		.USE_ADDRESS                    (1),
		.USE_WAITREQUEST                (0),
		.USE_WRITEBYTEENABLE            (0),
		.USE_OUTPUTENABLE               (0),
		.USE_RESETREQUEST               (0),
		.USE_IRQ                        (0),
		.USE_RESET_OUTPUT               (0),
		.ACTIVE_LOW_READ                (1),
		.ACTIVE_LOW_LOCK                (0),
		.ACTIVE_LOW_WRITE               (1),
		.ACTIVE_LOW_CHIPSELECT          (1),
		.ACTIVE_LOW_BYTEENABLE          (0),
		.ACTIVE_LOW_OUTPUTENABLE        (0),
		.ACTIVE_LOW_WRITEBYTEENABLE     (0),
		.ACTIVE_LOW_WAITREQUEST         (0),
		.ACTIVE_LOW_BEGINTRANSFER       (0),
		.CHIPSELECT_THROUGH_READLATENCY (0)
	) generic_tristate_controller_0 (
		.clk_clk              (altpll_0_c1_clk),                                                                //   clk.clk
		.reset_reset          (rst_controller_reset_out_reset),                                                 // reset.reset
		.uas_address          (generic_tristate_controller_0_uas_translator_avalon_anti_slave_0_address),       //   uas.address
		.uas_burstcount       (generic_tristate_controller_0_uas_translator_avalon_anti_slave_0_burstcount),    //      .burstcount
		.uas_read             (generic_tristate_controller_0_uas_translator_avalon_anti_slave_0_read),          //      .read
		.uas_write            (generic_tristate_controller_0_uas_translator_avalon_anti_slave_0_write),         //      .write
		.uas_waitrequest      (generic_tristate_controller_0_uas_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.uas_readdatavalid    (generic_tristate_controller_0_uas_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.uas_byteenable       (generic_tristate_controller_0_uas_translator_avalon_anti_slave_0_byteenable),    //      .byteenable
		.uas_readdata         (generic_tristate_controller_0_uas_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.uas_writedata        (generic_tristate_controller_0_uas_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.uas_lock             (generic_tristate_controller_0_uas_translator_avalon_anti_slave_0_lock),          //      .lock
		.uas_debugaccess      (generic_tristate_controller_0_uas_translator_avalon_anti_slave_0_debugaccess),   //      .debugaccess
		.tcm_write_n_out      (generic_tristate_controller_0_tcm_write_n_out),                                  //   tcm.write_n_out
		.tcm_read_n_out       (generic_tristate_controller_0_tcm_read_n_out),                                   //      .read_n_out
		.tcm_chipselect_n_out (generic_tristate_controller_0_tcm_chipselect_n_out),                             //      .chipselect_n_out
		.tcm_request          (generic_tristate_controller_0_tcm_request),                                      //      .request
		.tcm_grant            (generic_tristate_controller_0_tcm_grant),                                        //      .grant
		.tcm_address_out      (generic_tristate_controller_0_tcm_address_out),                                  //      .address_out
		.tcm_data_out         (generic_tristate_controller_0_tcm_data_out),                                     //      .data_out
		.tcm_data_outen       (generic_tristate_controller_0_tcm_data_outen),                                   //      .data_outen
		.tcm_data_in          (generic_tristate_controller_0_tcm_data_in)                                       //      .data_in
	);

	niosII_system_tristate_conduit_bridge_0 tristate_conduit_bridge_0 (
		.clk                                                    (altpll_0_c1_clk),                                                                          //   clk.clk
		.reset                                                  (rst_controller_reset_out_reset),                                                           // reset.reset
		.request                                                (tristate_conduit_pin_sharer_0_tcm_request),                                                //   tcs.request
		.grant                                                  (tristate_conduit_pin_sharer_0_tcm_grant),                                                  //      .grant
		.tcs_generic_tristate_controller_0_tcm_read_n_out       (tristate_conduit_pin_sharer_0_tcm_generic_tristate_controller_0_tcm_read_n_out_out),       //      .generic_tristate_controller_0_tcm_read_n_out_out
		.tcs_generic_tristate_controller_0_tcm_data_out         (tristate_conduit_pin_sharer_0_tcm_generic_tristate_controller_0_tcm_data_out_out),         //      .generic_tristate_controller_0_tcm_data_out_out
		.tcs_generic_tristate_controller_0_tcm_data_outen       (tristate_conduit_pin_sharer_0_tcm_generic_tristate_controller_0_tcm_data_out_outen),       //      .generic_tristate_controller_0_tcm_data_out_outen
		.tcs_generic_tristate_controller_0_tcm_data_in          (tristate_conduit_pin_sharer_0_tcm_generic_tristate_controller_0_tcm_data_out_in),          //      .generic_tristate_controller_0_tcm_data_out_in
		.tcs_generic_tristate_controller_0_tcm_chipselect_n_out (tristate_conduit_pin_sharer_0_tcm_generic_tristate_controller_0_tcm_chipselect_n_out_out), //      .generic_tristate_controller_0_tcm_chipselect_n_out_out
		.tcs_generic_tristate_controller_0_tcm_write_n_out      (tristate_conduit_pin_sharer_0_tcm_generic_tristate_controller_0_tcm_write_n_out_out),      //      .generic_tristate_controller_0_tcm_write_n_out_out
		.tcs_generic_tristate_controller_0_tcm_address_out      (tristate_conduit_pin_sharer_0_tcm_generic_tristate_controller_0_tcm_address_out_out),      //      .generic_tristate_controller_0_tcm_address_out_out
		.generic_tristate_controller_0_tcm_read_n_out           (tristate_conduit_bridge_0_out_generic_tristate_controller_0_tcm_read_n_out),               //   out.generic_tristate_controller_0_tcm_read_n_out
		.generic_tristate_controller_0_tcm_data_out             (tristate_conduit_bridge_0_out_generic_tristate_controller_0_tcm_data_out),                 //      .generic_tristate_controller_0_tcm_data_out
		.generic_tristate_controller_0_tcm_chipselect_n_out     (tristate_conduit_bridge_0_out_generic_tristate_controller_0_tcm_chipselect_n_out),         //      .generic_tristate_controller_0_tcm_chipselect_n_out
		.generic_tristate_controller_0_tcm_write_n_out          (tristate_conduit_bridge_0_out_generic_tristate_controller_0_tcm_write_n_out),              //      .generic_tristate_controller_0_tcm_write_n_out
		.generic_tristate_controller_0_tcm_address_out          (tristate_conduit_bridge_0_out_generic_tristate_controller_0_tcm_address_out)               //      .generic_tristate_controller_0_tcm_address_out
	);

	niosII_system_tristate_conduit_pin_sharer_0 tristate_conduit_pin_sharer_0 (
		.clk_clk                                            (altpll_0_c1_clk),                                                                          //   clk.clk
		.reset_reset                                        (rst_controller_reset_out_reset),                                                           // reset.reset
		.request                                            (tristate_conduit_pin_sharer_0_tcm_request),                                                //   tcm.request
		.grant                                              (tristate_conduit_pin_sharer_0_tcm_grant),                                                  //      .grant
		.generic_tristate_controller_0_tcm_address_out      (tristate_conduit_pin_sharer_0_tcm_generic_tristate_controller_0_tcm_address_out_out),      //      .generic_tristate_controller_0_tcm_address_out_out
		.generic_tristate_controller_0_tcm_read_n_out       (tristate_conduit_pin_sharer_0_tcm_generic_tristate_controller_0_tcm_read_n_out_out),       //      .generic_tristate_controller_0_tcm_read_n_out_out
		.generic_tristate_controller_0_tcm_write_n_out      (tristate_conduit_pin_sharer_0_tcm_generic_tristate_controller_0_tcm_write_n_out_out),      //      .generic_tristate_controller_0_tcm_write_n_out_out
		.generic_tristate_controller_0_tcm_data_out         (tristate_conduit_pin_sharer_0_tcm_generic_tristate_controller_0_tcm_data_out_out),         //      .generic_tristate_controller_0_tcm_data_out_out
		.generic_tristate_controller_0_tcm_data_in          (tristate_conduit_pin_sharer_0_tcm_generic_tristate_controller_0_tcm_data_out_in),          //      .generic_tristate_controller_0_tcm_data_out_in
		.generic_tristate_controller_0_tcm_data_outen       (tristate_conduit_pin_sharer_0_tcm_generic_tristate_controller_0_tcm_data_out_outen),       //      .generic_tristate_controller_0_tcm_data_out_outen
		.generic_tristate_controller_0_tcm_chipselect_n_out (tristate_conduit_pin_sharer_0_tcm_generic_tristate_controller_0_tcm_chipselect_n_out_out), //      .generic_tristate_controller_0_tcm_chipselect_n_out_out
		.tcs0_request                                       (generic_tristate_controller_0_tcm_request),                                                //  tcs0.request
		.tcs0_grant                                         (generic_tristate_controller_0_tcm_grant),                                                  //      .grant
		.tcs0_address_out                                   (generic_tristate_controller_0_tcm_address_out),                                            //      .address_out
		.tcs0_read_n_out                                    (generic_tristate_controller_0_tcm_read_n_out),                                             //      .read_n_out
		.tcs0_write_n_out                                   (generic_tristate_controller_0_tcm_write_n_out),                                            //      .write_n_out
		.tcs0_data_out                                      (generic_tristate_controller_0_tcm_data_out),                                               //      .data_out
		.tcs0_data_in                                       (generic_tristate_controller_0_tcm_data_in),                                                //      .data_in
		.tcs0_data_outen                                    (generic_tristate_controller_0_tcm_data_outen),                                             //      .data_outen
		.tcs0_chipselect_n_out                              (generic_tristate_controller_0_tcm_chipselect_n_out)                                        //      .chipselect_n_out
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (25),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (25),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_qsys_0_instruction_master_translator (
		.clk                   (altpll_0_c1_clk),                                                                    //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                     //                     reset.reset
		.uav_address           (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (nios2_qsys_0_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (nios2_qsys_0_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read               (nios2_qsys_0_instruction_master_read),                                               //                          .read
		.av_readdata           (nios2_qsys_0_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (nios2_qsys_0_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                               //               (terminated)
		.av_byteenable         (4'b1111),                                                                            //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                               //               (terminated)
		.av_begintransfer      (1'b0),                                                                               //               (terminated)
		.av_chipselect         (1'b0),                                                                               //               (terminated)
		.av_write              (1'b0),                                                                               //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                               //               (terminated)
		.av_lock               (1'b0),                                                                               //               (terminated)
		.av_debugaccess        (1'b0),                                                                               //               (terminated)
		.uav_clken             (),                                                                                   //               (terminated)
		.av_clken              (1'b1)                                                                                //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (25),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (25),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_qsys_0_data_master_translator (
		.clk                   (altpll_0_c1_clk),                                                             //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                              //                     reset.reset
		.uav_address           (nios2_qsys_0_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (nios2_qsys_0_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (nios2_qsys_0_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (nios2_qsys_0_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (nios2_qsys_0_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (nios2_qsys_0_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (nios2_qsys_0_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (nios2_qsys_0_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (nios2_qsys_0_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (nios2_qsys_0_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (nios2_qsys_0_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (nios2_qsys_0_data_master_byteenable),                                         //                          .byteenable
		.av_read               (nios2_qsys_0_data_master_read),                                               //                          .read
		.av_readdata           (nios2_qsys_0_data_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (nios2_qsys_0_data_master_readdatavalid),                                      //                          .readdatavalid
		.av_write              (nios2_qsys_0_data_master_write),                                              //                          .write
		.av_writedata          (nios2_qsys_0_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (nios2_qsys_0_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount         (1'b1),                                                                        //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                        //               (terminated)
		.av_begintransfer      (1'b0),                                                                        //               (terminated)
		.av_chipselect         (1'b0),                                                                        //               (terminated)
		.av_lock               (1'b0),                                                                        //               (terminated)
		.uav_clken             (),                                                                            //               (terminated)
		.av_clken              (1'b1)                                                                         //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) nios2_qsys_0_jtag_debug_module_translator (
		.clk                   (altpll_0_c1_clk),                                                                           //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                            //                    reset.reset
		.uav_address           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                          //              (terminated)
		.av_beginbursttransfer (),                                                                                          //              (terminated)
		.av_burstcount         (),                                                                                          //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                      //              (terminated)
		.av_waitrequest        (1'b0),                                                                                      //              (terminated)
		.av_writebyteenable    (),                                                                                          //              (terminated)
		.av_lock               (),                                                                                          //              (terminated)
		.av_clken              (),                                                                                          //              (terminated)
		.uav_clken             (1'b0),                                                                                      //              (terminated)
		.av_outputenable       ()                                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (12),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) onchip_memory2_0_s1_translator (
		.clk                   (altpll_0_c1_clk),                                                                //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                 //                    reset.reset
		.uav_address           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (onchip_memory2_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (onchip_memory2_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                               //              (terminated)
		.av_begintransfer      (),                                                                               //              (terminated)
		.av_beginbursttransfer (),                                                                               //              (terminated)
		.av_burstcount         (),                                                                               //              (terminated)
		.av_readdatavalid      (1'b0),                                                                           //              (terminated)
		.av_waitrequest        (1'b0),                                                                           //              (terminated)
		.av_writebyteenable    (),                                                                               //              (terminated)
		.av_lock               (),                                                                               //              (terminated)
		.uav_clken             (1'b0),                                                                           //              (terminated)
		.av_debugaccess        (),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (22),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sdram_0_s1_translator (
		.clk                   (altpll_0_c1_clk),                                                       //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address           (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sdram_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sdram_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sdram_0_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sdram_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sdram_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (sdram_0_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (sdram_0_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (sdram_0_s1_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (sdram_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (18),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sram_0_avalon_sram_slave_translator (
		.clk                   (altpll_0_c1_clk),                                                                     //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                      //                    reset.reset
		.uav_address           (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_begintransfer      (),                                                                                    //              (terminated)
		.av_beginbursttransfer (),                                                                                    //              (terminated)
		.av_burstcount         (),                                                                                    //              (terminated)
		.av_waitrequest        (1'b0),                                                                                //              (terminated)
		.av_writebyteenable    (),                                                                                    //              (terminated)
		.av_lock               (),                                                                                    //              (terminated)
		.av_chipselect         (),                                                                                    //              (terminated)
		.av_clken              (),                                                                                    //              (terminated)
		.uav_clken             (1'b0),                                                                                //              (terminated)
		.av_debugaccess        (),                                                                                    //              (terminated)
		.av_outputenable       ()                                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sd_card_spi_master_spi_control_port_translator (
		.clk                   (altpll_0_c1_clk),                                                                                //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                                 //                    reset.reset
		.uav_address           (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sd_card_spi_master_spi_control_port_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sd_card_spi_master_spi_control_port_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sd_card_spi_master_spi_control_port_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sd_card_spi_master_spi_control_port_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sd_card_spi_master_spi_control_port_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (sd_card_spi_master_spi_control_port_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                               //              (terminated)
		.av_beginbursttransfer (),                                                                                               //              (terminated)
		.av_burstcount         (),                                                                                               //              (terminated)
		.av_byteenable         (),                                                                                               //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                           //              (terminated)
		.av_waitrequest        (1'b0),                                                                                           //              (terminated)
		.av_writebyteenable    (),                                                                                               //              (terminated)
		.av_lock               (),                                                                                               //              (terminated)
		.av_clken              (),                                                                                               //              (terminated)
		.uav_clken             (1'b0),                                                                                           //              (terminated)
		.av_debugaccess        (),                                                                                               //              (terminated)
		.av_outputenable       ()                                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (22),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (1),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) generic_tristate_controller_0_uas_translator (
		.clk                   (altpll_0_c1_clk),                                                                              //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                               //                    reset.reset
		.uav_address           (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (generic_tristate_controller_0_uas_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (generic_tristate_controller_0_uas_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (generic_tristate_controller_0_uas_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (generic_tristate_controller_0_uas_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (generic_tristate_controller_0_uas_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount         (generic_tristate_controller_0_uas_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable         (generic_tristate_controller_0_uas_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (generic_tristate_controller_0_uas_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (generic_tristate_controller_0_uas_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_lock               (generic_tristate_controller_0_uas_translator_avalon_anti_slave_0_lock),                        //                         .lock
		.av_debugaccess        (generic_tristate_controller_0_uas_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer      (),                                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                                             //              (terminated)
		.av_writebyteenable    (),                                                                                             //              (terminated)
		.av_chipselect         (),                                                                                             //              (terminated)
		.av_clken              (),                                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                                         //              (terminated)
		.av_outputenable       ()                                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) altpll_0_pll_slave_translator (
		.clk                   (clk_clk),                                                                       //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                            //                    reset.reset
		.uav_address           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (altpll_0_pll_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (altpll_0_pll_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (altpll_0_pll_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (altpll_0_pll_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (altpll_0_pll_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_waitrequest        (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sysid_qsys_0_control_slave_translator (
		.clk                   (altpll_0_c1_clk),                                                                       //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                        //                    reset.reset
		.uav_address           (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata           (sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write              (),                                                                                      //              (terminated)
		.av_read               (),                                                                                      //              (terminated)
		.av_writedata          (),                                                                                      //              (terminated)
		.av_begintransfer      (),                                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                                      //              (terminated)
		.av_burstcount         (),                                                                                      //              (terminated)
		.av_byteenable         (),                                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                                      //              (terminated)
		.av_lock               (),                                                                                      //              (terminated)
		.av_chipselect         (),                                                                                      //              (terminated)
		.av_clken              (),                                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                                  //              (terminated)
		.av_debugaccess        (),                                                                                      //              (terminated)
		.av_outputenable       ()                                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_0_s1_translator (
		.clk                   (altpll_0_c1_clk),                                                       //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (timer_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (timer_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (timer_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (timer_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (timer_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_0_avalon_jtag_slave_translator (
		.clk                   (altpll_0_c1_clk),                                                                          //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                           //                    reset.reset
		.uav_address           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                                         //              (terminated)
		.av_burstcount         (),                                                                                         //              (terminated)
		.av_byteenable         (),                                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                                         //              (terminated)
		.av_lock               (),                                                                                         //              (terminated)
		.av_clken              (),                                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                                     //              (terminated)
		.av_debugaccess        (),                                                                                         //              (terminated)
		.av_outputenable       ()                                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) character_lcd_0_avalon_lcd_slave_translator (
		.clk                   (altpll_0_c1_clk),                                                                             //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                              //                    reset.reset
		.uav_address           (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                            //              (terminated)
		.av_beginbursttransfer (),                                                                                            //              (terminated)
		.av_burstcount         (),                                                                                            //              (terminated)
		.av_byteenable         (),                                                                                            //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                        //              (terminated)
		.av_writebyteenable    (),                                                                                            //              (terminated)
		.av_lock               (),                                                                                            //              (terminated)
		.av_clken              (),                                                                                            //              (terminated)
		.uav_clken             (1'b0),                                                                                        //              (terminated)
		.av_debugaccess        (),                                                                                            //              (terminated)
		.av_outputenable       ()                                                                                             //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) green_leds_s1_translator (
		.clk                   (altpll_0_c1_clk),                                                          //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                           //                    reset.reset
		.uav_address           (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (green_leds_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (green_leds_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (green_leds_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (green_leds_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (green_leds_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                         //              (terminated)
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_byteenable         (),                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.av_clken              (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) switch_s1_translator (
		.clk                   (altpll_0_c1_clk),                                                      //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                       //                    reset.reset
		.uav_address           (switch_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (switch_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (switch_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (switch_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (switch_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (switch_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (switch_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (switch_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (switch_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (switch_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (switch_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (switch_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata           (switch_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write              (),                                                                     //              (terminated)
		.av_read               (),                                                                     //              (terminated)
		.av_writedata          (),                                                                     //              (terminated)
		.av_begintransfer      (),                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                     //              (terminated)
		.av_burstcount         (),                                                                     //              (terminated)
		.av_byteenable         (),                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                 //              (terminated)
		.av_waitrequest        (1'b0),                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                     //              (terminated)
		.av_lock               (),                                                                     //              (terminated)
		.av_chipselect         (),                                                                     //              (terminated)
		.av_clken              (),                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                 //              (terminated)
		.av_debugaccess        (),                                                                     //              (terminated)
		.av_outputenable       ()                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) audio_0_avalon_audio_slave_translator (
		.clk                   (up_clocks_1_audio_clk_clk),                                                             //                      clk.clk
		.reset                 (rst_controller_002_reset_out_reset),                                                    //                    reset.reset
		.uav_address           (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (audio_0_avalon_audio_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (audio_0_avalon_audio_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (audio_0_avalon_audio_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (audio_0_avalon_audio_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (audio_0_avalon_audio_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (audio_0_avalon_audio_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                                      //              (terminated)
		.av_burstcount         (),                                                                                      //              (terminated)
		.av_byteenable         (),                                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                                      //              (terminated)
		.av_lock               (),                                                                                      //              (terminated)
		.av_clken              (),                                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                                  //              (terminated)
		.av_debugaccess        (),                                                                                      //              (terminated)
		.av_outputenable       ()                                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) audio_and_video_config_0_avalon_av_config_slave_translator (
		.clk                   (up_clocks_1_audio_clk_clk),                                                                                  //                      clk.clk
		.reset                 (rst_controller_002_reset_out_reset),                                                                         //                    reset.reset
		.uav_address           (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_begintransfer      (),                                                                                                           //              (terminated)
		.av_beginbursttransfer (),                                                                                                           //              (terminated)
		.av_burstcount         (),                                                                                                           //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                                       //              (terminated)
		.av_writebyteenable    (),                                                                                                           //              (terminated)
		.av_lock               (),                                                                                                           //              (terminated)
		.av_chipselect         (),                                                                                                           //              (terminated)
		.av_clken              (),                                                                                                           //              (terminated)
		.uav_clken             (1'b0),                                                                                                       //              (terminated)
		.av_debugaccess        (),                                                                                                           //              (terminated)
		.av_outputenable       ()                                                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) i2c_scl_s1_translator (
		.clk                   (altpll_0_c1_clk),                                                       //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address           (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (i2c_scl_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (i2c_scl_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (i2c_scl_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (i2c_scl_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (i2c_scl_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) i2c_sda_s1_translator (
		.clk                   (altpll_0_c1_clk),                                                       //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address           (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (i2c_sda_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (i2c_sda_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (i2c_sda_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (i2c_sda_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (i2c_sda_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) i2c_scl_2_s1_translator (
		.clk                   (altpll_0_c1_clk),                                                         //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                          //                    reset.reset
		.uav_address           (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (i2c_scl_2_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (i2c_scl_2_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (i2c_scl_2_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (i2c_scl_2_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (i2c_scl_2_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                        //              (terminated)
		.av_begintransfer      (),                                                                        //              (terminated)
		.av_beginbursttransfer (),                                                                        //              (terminated)
		.av_burstcount         (),                                                                        //              (terminated)
		.av_byteenable         (),                                                                        //              (terminated)
		.av_readdatavalid      (1'b0),                                                                    //              (terminated)
		.av_waitrequest        (1'b0),                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                        //              (terminated)
		.av_lock               (),                                                                        //              (terminated)
		.av_clken              (),                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                    //              (terminated)
		.av_debugaccess        (),                                                                        //              (terminated)
		.av_outputenable       ()                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) i2c_sda_2_s1_translator (
		.clk                   (altpll_0_c1_clk),                                                         //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                          //                    reset.reset
		.uav_address           (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (i2c_sda_2_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (i2c_sda_2_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (i2c_sda_2_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (i2c_sda_2_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (i2c_sda_2_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                        //              (terminated)
		.av_begintransfer      (),                                                                        //              (terminated)
		.av_beginbursttransfer (),                                                                        //              (terminated)
		.av_burstcount         (),                                                                        //              (terminated)
		.av_byteenable         (),                                                                        //              (terminated)
		.av_readdatavalid      (1'b0),                                                                    //              (terminated)
		.av_waitrequest        (1'b0),                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                        //              (terminated)
		.av_lock               (),                                                                        //              (terminated)
		.av_clken              (),                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                    //              (terminated)
		.av_debugaccess        (),                                                                        //              (terminated)
		.av_outputenable       ()                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) drum_out_s1_translator (
		.clk                   (altpll_0_c1_clk),                                                        //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                         //                    reset.reset
		.uav_address           (drum_out_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (drum_out_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (drum_out_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (drum_out_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (drum_out_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (drum_out_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (drum_out_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (drum_out_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (drum_out_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (drum_out_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (drum_out_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (drum_out_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (drum_out_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (drum_out_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (drum_out_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (drum_out_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                       //              (terminated)
		.av_begintransfer      (),                                                                       //              (terminated)
		.av_beginbursttransfer (),                                                                       //              (terminated)
		.av_burstcount         (),                                                                       //              (terminated)
		.av_byteenable         (),                                                                       //              (terminated)
		.av_readdatavalid      (1'b0),                                                                   //              (terminated)
		.av_waitrequest        (1'b0),                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                       //              (terminated)
		.av_lock               (),                                                                       //              (terminated)
		.av_clken              (),                                                                       //              (terminated)
		.uav_clken             (1'b0),                                                                   //              (terminated)
		.av_debugaccess        (),                                                                       //              (terminated)
		.av_outputenable       ()                                                                        //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (95),
		.PKT_PROTECTION_L          (93),
		.PKT_BEGIN_BURST           (80),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.PKT_BURST_TYPE_H          (77),
		.PKT_BURST_TYPE_L          (76),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_TRANS_EXCLUSIVE       (66),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (87),
		.PKT_THREAD_ID_H           (92),
		.PKT_THREAD_ID_L           (92),
		.PKT_CACHE_H               (99),
		.PKT_CACHE_L               (96),
		.PKT_DATA_SIDEBAND_H       (79),
		.PKT_DATA_SIDEBAND_L       (79),
		.PKT_QOS_H                 (81),
		.PKT_QOS_L                 (81),
		.PKT_ADDR_SIDEBAND_H       (78),
		.PKT_ADDR_SIDEBAND_L       (78),
		.ST_DATA_W                 (102),
		.ST_CHANNEL_W              (20),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (4'b0000)
	) nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (altpll_0_c1_clk),                                                                             //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.av_address       (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_rsp_src_valid),                                                                       //        rp.valid
		.rp_data          (limiter_rsp_src_data),                                                                        //          .data
		.rp_channel       (limiter_rsp_src_channel),                                                                     //          .channel
		.rp_startofpacket (limiter_rsp_src_startofpacket),                                                               //          .startofpacket
		.rp_endofpacket   (limiter_rsp_src_endofpacket),                                                                 //          .endofpacket
		.rp_ready         (limiter_rsp_src_ready)                                                                        //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (95),
		.PKT_PROTECTION_L          (93),
		.PKT_BEGIN_BURST           (80),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.PKT_BURST_TYPE_H          (77),
		.PKT_BURST_TYPE_L          (76),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_TRANS_EXCLUSIVE       (66),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (87),
		.PKT_THREAD_ID_H           (92),
		.PKT_THREAD_ID_L           (92),
		.PKT_CACHE_H               (99),
		.PKT_CACHE_L               (96),
		.PKT_DATA_SIDEBAND_H       (79),
		.PKT_DATA_SIDEBAND_L       (79),
		.PKT_QOS_H                 (81),
		.PKT_QOS_L                 (81),
		.PKT_ADDR_SIDEBAND_H       (78),
		.PKT_ADDR_SIDEBAND_L       (78),
		.ST_DATA_W                 (102),
		.ST_CHANNEL_W              (20),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent (
		.clk              (altpll_0_c1_clk),                                                                      //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.av_address       (nios2_qsys_0_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (nios2_qsys_0_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (nios2_qsys_0_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (nios2_qsys_0_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (nios2_qsys_0_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (nios2_qsys_0_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (nios2_qsys_0_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_001_rsp_src_valid),                                                            //        rp.valid
		.rp_data          (limiter_001_rsp_src_data),                                                             //          .data
		.rp_channel       (limiter_001_rsp_src_channel),                                                          //          .channel
		.rp_startofpacket (limiter_001_rsp_src_startofpacket),                                                    //          .startofpacket
		.rp_endofpacket   (limiter_001_rsp_src_endofpacket),                                                      //          .endofpacket
		.rp_ready         (limiter_001_rsp_src_ready)                                                             //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (80),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (87),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (95),
		.PKT_PROTECTION_L          (93),
		.PKT_RESPONSE_STATUS_H     (101),
		.PKT_RESPONSE_STATUS_L     (100),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.ST_CHANNEL_W              (20),
		.ST_DATA_W                 (102),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c1_clk),                                                                                     //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                      //       clk_reset.reset
		.m0_address              (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                              //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                              //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                               //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                            //                .channel
		.rf_sink_ready           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (103),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c1_clk),                                                                                     //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                      // clk_reset.reset
		.in_data           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                                // (terminated)
		.csr_readdata      (),                                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                // (terminated)
		.almost_full_data  (),                                                                                                    // (terminated)
		.almost_empty_data (),                                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                                // (terminated)
		.out_empty         (),                                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                                // (terminated)
		.out_error         (),                                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                                // (terminated)
		.out_channel       ()                                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (80),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (87),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (95),
		.PKT_PROTECTION_L          (93),
		.PKT_RESPONSE_STATUS_H     (101),
		.PKT_RESPONSE_STATUS_L     (100),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.ST_CHANNEL_W              (20),
		.ST_DATA_W                 (102),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c1_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_001_src_ready),                                                               //              cp.ready
		.cp_valid                (cmd_xbar_mux_001_src_valid),                                                               //                .valid
		.cp_data                 (cmd_xbar_mux_001_src_data),                                                                //                .data
		.cp_startofpacket        (cmd_xbar_mux_001_src_startofpacket),                                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_001_src_endofpacket),                                                         //                .endofpacket
		.cp_channel              (cmd_xbar_mux_001_src_channel),                                                             //                .channel
		.rf_sink_ready           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (103),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c1_clk),                                                                          //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (62),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (42),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (43),
		.PKT_TRANS_POSTED          (44),
		.PKT_TRANS_WRITE           (45),
		.PKT_TRANS_READ            (46),
		.PKT_TRANS_LOCK            (47),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (64),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (54),
		.PKT_BURSTWRAP_L           (52),
		.PKT_BYTE_CNT_H            (51),
		.PKT_BYTE_CNT_L            (49),
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_RESPONSE_STATUS_H     (83),
		.PKT_RESPONSE_STATUS_L     (82),
		.PKT_BURST_SIZE_H          (57),
		.PKT_BURST_SIZE_L          (55),
		.ST_CHANNEL_W              (20),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sdram_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c1_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                     //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                     //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                      //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                               //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                   //                .channel
		.rf_sink_ready           (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c1_clk),                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (62),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (42),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (43),
		.PKT_TRANS_POSTED          (44),
		.PKT_TRANS_WRITE           (45),
		.PKT_TRANS_READ            (46),
		.PKT_TRANS_LOCK            (47),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (64),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (54),
		.PKT_BURSTWRAP_L           (52),
		.PKT_BYTE_CNT_H            (51),
		.PKT_BYTE_CNT_L            (49),
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_RESPONSE_STATUS_H     (83),
		.PKT_RESPONSE_STATUS_L     (82),
		.PKT_BURST_SIZE_H          (57),
		.PKT_BURST_SIZE_L          (55),
		.ST_CHANNEL_W              (20),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c1_clk),                                                                               //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                //       clk_reset.reset
		.m0_address              (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_001_source0_ready),                                                               //              cp.ready
		.cp_valid                (burst_adapter_001_source0_valid),                                                               //                .valid
		.cp_data                 (burst_adapter_001_source0_data),                                                                //                .data
		.cp_startofpacket        (burst_adapter_001_source0_startofpacket),                                                       //                .startofpacket
		.cp_endofpacket          (burst_adapter_001_source0_endofpacket),                                                         //                .endofpacket
		.cp_channel              (burst_adapter_001_source0_channel),                                                             //                .channel
		.rf_sink_ready           (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (3),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c1_clk),                                                                               //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                // clk_reset.reset
		.in_data           (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                          // (terminated)
		.csr_readdata      (),                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                          // (terminated)
		.almost_full_data  (),                                                                                              // (terminated)
		.almost_empty_data (),                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                          // (terminated)
		.out_empty         (),                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                          // (terminated)
		.out_error         (),                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                          // (terminated)
		.out_channel       ()                                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (80),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (87),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (95),
		.PKT_PROTECTION_L          (93),
		.PKT_RESPONSE_STATUS_H     (101),
		.PKT_RESPONSE_STATUS_L     (100),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.ST_CHANNEL_W              (20),
		.ST_DATA_W                 (102),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c1_clk),                                                                                          //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                           //       clk_reset.reset
		.m0_address              (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_004_src_ready),                                                                               //              cp.ready
		.cp_valid                (cmd_xbar_mux_004_src_valid),                                                                               //                .valid
		.cp_data                 (cmd_xbar_mux_004_src_data),                                                                                //                .data
		.cp_startofpacket        (cmd_xbar_mux_004_src_startofpacket),                                                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_004_src_endofpacket),                                                                         //                .endofpacket
		.cp_channel              (cmd_xbar_mux_004_src_channel),                                                                             //                .channel
		.rf_sink_ready           (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (103),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c1_clk),                                                                                          //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                           // clk_reset.reset
		.in_data           (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                                     // (terminated)
		.csr_readdata      (),                                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                     // (terminated)
		.almost_full_data  (),                                                                                                         // (terminated)
		.almost_empty_data (),                                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                                     // (terminated)
		.out_empty         (),                                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                                     // (terminated)
		.out_error         (),                                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                                     // (terminated)
		.out_channel       ()                                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (53),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (33),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (34),
		.PKT_TRANS_POSTED          (35),
		.PKT_TRANS_WRITE           (36),
		.PKT_TRANS_READ            (37),
		.PKT_TRANS_LOCK            (38),
		.PKT_SRC_ID_H              (59),
		.PKT_SRC_ID_L              (55),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (60),
		.PKT_BURSTWRAP_H           (45),
		.PKT_BURSTWRAP_L           (43),
		.PKT_BYTE_CNT_H            (42),
		.PKT_BYTE_CNT_L            (40),
		.PKT_PROTECTION_H          (68),
		.PKT_PROTECTION_L          (66),
		.PKT_RESPONSE_STATUS_H     (74),
		.PKT_RESPONSE_STATUS_L     (73),
		.PKT_BURST_SIZE_H          (48),
		.PKT_BURST_SIZE_L          (46),
		.ST_CHANNEL_W              (20),
		.ST_DATA_W                 (75),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c1_clk),                                                                                        //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                         //       clk_reset.reset
		.m0_address              (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_002_source0_ready),                                                                        //              cp.ready
		.cp_valid                (burst_adapter_002_source0_valid),                                                                        //                .valid
		.cp_data                 (burst_adapter_002_source0_data),                                                                         //                .data
		.cp_startofpacket        (burst_adapter_002_source0_startofpacket),                                                                //                .startofpacket
		.cp_endofpacket          (burst_adapter_002_source0_endofpacket),                                                                  //                .endofpacket
		.cp_channel              (burst_adapter_002_source0_channel),                                                                      //                .channel
		.rf_sink_ready           (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (76),
		.FIFO_DEPTH          (4),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c1_clk),                                                                                        //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                         // clk_reset.reset
		.in_data           (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                                   // (terminated)
		.csr_readdata      (),                                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                   // (terminated)
		.almost_full_data  (),                                                                                                       // (terminated)
		.almost_empty_data (),                                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                                   // (terminated)
		.out_empty         (),                                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                                   // (terminated)
		.out_error         (),                                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                                   // (terminated)
		.out_channel       ()                                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (80),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (87),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (95),
		.PKT_PROTECTION_L          (93),
		.PKT_RESPONSE_STATUS_H     (101),
		.PKT_RESPONSE_STATUS_L     (100),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.ST_CHANNEL_W              (20),
		.ST_DATA_W                 (102),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) altpll_0_pll_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                 //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                      //       clk_reset.reset
		.m0_address              (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_out_ready),                                                                       //              cp.ready
		.cp_valid                (crosser_out_valid),                                                                       //                .valid
		.cp_data                 (crosser_out_data),                                                                        //                .data
		.cp_startofpacket        (crosser_out_startofpacket),                                                               //                .startofpacket
		.cp_endofpacket          (crosser_out_endofpacket),                                                                 //                .endofpacket
		.cp_channel              (crosser_out_channel),                                                                     //                .channel
		.rf_sink_ready           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (103),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                 //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                      // clk_reset.reset
		.in_data           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_startofpacket  (1'b0),                                                                              // (terminated)
		.in_endofpacket    (1'b0),                                                                              // (terminated)
		.out_startofpacket (),                                                                                  // (terminated)
		.out_endofpacket   (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (80),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (87),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (95),
		.PKT_PROTECTION_L          (93),
		.PKT_RESPONSE_STATUS_H     (101),
		.PKT_RESPONSE_STATUS_L     (100),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.ST_CHANNEL_W              (20),
		.ST_DATA_W                 (102),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c1_clk),                                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                  //       clk_reset.reset
		.m0_address              (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src7_ready),                                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src7_valid),                                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src7_data),                                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src7_startofpacket),                                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src7_endofpacket),                                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src7_channel),                                                                 //                .channel
		.rf_sink_ready           (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (103),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c1_clk),                                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                  // clk_reset.reset
		.in_data           (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                           // (terminated)
		.csr_read          (1'b0),                                                                                            // (terminated)
		.csr_write         (1'b0),                                                                                            // (terminated)
		.csr_readdata      (),                                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                            // (terminated)
		.almost_full_data  (),                                                                                                // (terminated)
		.almost_empty_data (),                                                                                                // (terminated)
		.in_empty          (1'b0),                                                                                            // (terminated)
		.out_empty         (),                                                                                                // (terminated)
		.in_error          (1'b0),                                                                                            // (terminated)
		.out_error         (),                                                                                                // (terminated)
		.in_channel        (1'b0),                                                                                            // (terminated)
		.out_channel       ()                                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (80),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (87),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (95),
		.PKT_PROTECTION_L          (93),
		.PKT_RESPONSE_STATUS_H     (101),
		.PKT_RESPONSE_STATUS_L     (100),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.ST_CHANNEL_W              (20),
		.ST_DATA_W                 (102),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) timer_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c1_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src8_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src8_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src8_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src8_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src8_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src8_channel),                                                 //                .channel
		.rf_sink_ready           (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (103),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c1_clk),                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (80),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (87),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (95),
		.PKT_PROTECTION_L          (93),
		.PKT_RESPONSE_STATUS_H     (101),
		.PKT_RESPONSE_STATUS_L     (100),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.ST_CHANNEL_W              (20),
		.ST_DATA_W                 (102),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c1_clk),                                                                                    //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                     //       clk_reset.reset
		.m0_address              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src9_ready),                                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src9_valid),                                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_001_src9_data),                                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src9_startofpacket),                                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src9_endofpacket),                                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src9_channel),                                                                    //                .channel
		.rf_sink_ready           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (103),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c1_clk),                                                                                    //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                     // clk_reset.reset
		.in_data           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (53),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (33),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (34),
		.PKT_TRANS_POSTED          (35),
		.PKT_TRANS_WRITE           (36),
		.PKT_TRANS_READ            (37),
		.PKT_TRANS_LOCK            (38),
		.PKT_SRC_ID_H              (59),
		.PKT_SRC_ID_L              (55),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (60),
		.PKT_BURSTWRAP_H           (45),
		.PKT_BURSTWRAP_L           (43),
		.PKT_BYTE_CNT_H            (42),
		.PKT_BYTE_CNT_L            (40),
		.PKT_PROTECTION_H          (68),
		.PKT_PROTECTION_L          (66),
		.PKT_RESPONSE_STATUS_H     (74),
		.PKT_RESPONSE_STATUS_L     (73),
		.PKT_BURST_SIZE_H          (48),
		.PKT_BURST_SIZE_L          (46),
		.ST_CHANNEL_W              (20),
		.ST_DATA_W                 (75),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c1_clk),                                                                                       //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                        //       clk_reset.reset
		.m0_address              (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_003_source0_ready),                                                                       //              cp.ready
		.cp_valid                (burst_adapter_003_source0_valid),                                                                       //                .valid
		.cp_data                 (burst_adapter_003_source0_data),                                                                        //                .data
		.cp_startofpacket        (burst_adapter_003_source0_startofpacket),                                                               //                .startofpacket
		.cp_endofpacket          (burst_adapter_003_source0_endofpacket),                                                                 //                .endofpacket
		.cp_channel              (burst_adapter_003_source0_channel),                                                                     //                .channel
		.rf_sink_ready           (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (76),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c1_clk),                                                                                       //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                        // clk_reset.reset
		.in_data           (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                                  // (terminated)
		.csr_readdata      (),                                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                  // (terminated)
		.almost_full_data  (),                                                                                                      // (terminated)
		.almost_empty_data (),                                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                                  // (terminated)
		.out_empty         (),                                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                                  // (terminated)
		.out_error         (),                                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                                  // (terminated)
		.out_channel       ()                                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (80),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (87),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (95),
		.PKT_PROTECTION_L          (93),
		.PKT_RESPONSE_STATUS_H     (101),
		.PKT_RESPONSE_STATUS_L     (100),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.ST_CHANNEL_W              (20),
		.ST_DATA_W                 (102),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) green_leds_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c1_clk),                                                                    //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src11_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src11_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src11_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src11_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src11_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src11_channel),                                                   //                .channel
		.rf_sink_ready           (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (103),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c1_clk),                                                                    //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (80),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (87),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (95),
		.PKT_PROTECTION_L          (93),
		.PKT_RESPONSE_STATUS_H     (101),
		.PKT_RESPONSE_STATUS_L     (100),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.ST_CHANNEL_W              (20),
		.ST_DATA_W                 (102),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) switch_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c1_clk),                                                                //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (switch_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (switch_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (switch_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (switch_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (switch_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (switch_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (switch_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (switch_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (switch_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (switch_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (switch_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (switch_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (switch_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (switch_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (switch_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (switch_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src12_ready),                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src12_valid),                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_001_src12_data),                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src12_startofpacket),                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src12_endofpacket),                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src12_channel),                                               //                .channel
		.rf_sink_ready           (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (103),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c1_clk),                                                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (80),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (87),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (95),
		.PKT_PROTECTION_L          (93),
		.PKT_RESPONSE_STATUS_H     (101),
		.PKT_RESPONSE_STATUS_L     (100),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.ST_CHANNEL_W              (20),
		.ST_DATA_W                 (102),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (up_clocks_1_audio_clk_clk),                                                                       //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                              //       clk_reset.reset
		.m0_address              (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_001_out_ready),                                                                           //              cp.ready
		.cp_valid                (crosser_001_out_valid),                                                                           //                .valid
		.cp_data                 (crosser_001_out_data),                                                                            //                .data
		.cp_startofpacket        (crosser_001_out_startofpacket),                                                                   //                .startofpacket
		.cp_endofpacket          (crosser_001_out_endofpacket),                                                                     //                .endofpacket
		.cp_channel              (crosser_001_out_channel),                                                                         //                .channel
		.rf_sink_ready           (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (103),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (up_clocks_1_audio_clk_clk),                                                                       //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                              // clk_reset.reset
		.in_data           (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                           // (terminated)
		.csr_read          (1'b0),                                                                                            // (terminated)
		.csr_write         (1'b0),                                                                                            // (terminated)
		.csr_readdata      (),                                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                            // (terminated)
		.almost_full_data  (),                                                                                                // (terminated)
		.almost_empty_data (),                                                                                                // (terminated)
		.in_empty          (1'b0),                                                                                            // (terminated)
		.out_empty         (),                                                                                                // (terminated)
		.in_error          (1'b0),                                                                                            // (terminated)
		.out_error         (),                                                                                                // (terminated)
		.in_channel        (1'b0),                                                                                            // (terminated)
		.out_channel       ()                                                                                                 // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (up_clocks_1_audio_clk_clk),                                                                 //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_startofpacket  (1'b0),                                                                                      // (terminated)
		.in_endofpacket    (1'b0),                                                                                      // (terminated)
		.out_startofpacket (),                                                                                          // (terminated)
		.out_endofpacket   (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (80),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (87),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (95),
		.PKT_PROTECTION_L          (93),
		.PKT_RESPONSE_STATUS_H     (101),
		.PKT_RESPONSE_STATUS_L     (100),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.ST_CHANNEL_W              (20),
		.ST_DATA_W                 (102),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (up_clocks_1_audio_clk_clk),                                                                                            //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                                                   //       clk_reset.reset
		.m0_address              (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_002_out_ready),                                                                                                //              cp.ready
		.cp_valid                (crosser_002_out_valid),                                                                                                //                .valid
		.cp_data                 (crosser_002_out_data),                                                                                                 //                .data
		.cp_startofpacket        (crosser_002_out_startofpacket),                                                                                        //                .startofpacket
		.cp_endofpacket          (crosser_002_out_endofpacket),                                                                                          //                .endofpacket
		.cp_channel              (crosser_002_out_channel),                                                                                              //                .channel
		.rf_sink_ready           (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (103),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (up_clocks_1_audio_clk_clk),                                                                                            //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                                                   // clk_reset.reset
		.in_data           (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                                // (terminated)
		.csr_read          (1'b0),                                                                                                                 // (terminated)
		.csr_write         (1'b0),                                                                                                                 // (terminated)
		.csr_readdata      (),                                                                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                                 // (terminated)
		.almost_full_data  (),                                                                                                                     // (terminated)
		.almost_empty_data (),                                                                                                                     // (terminated)
		.in_empty          (1'b0),                                                                                                                 // (terminated)
		.out_empty         (),                                                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                                                 // (terminated)
		.out_error         (),                                                                                                                     // (terminated)
		.in_channel        (1'b0),                                                                                                                 // (terminated)
		.out_channel       ()                                                                                                                      // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (up_clocks_1_audio_clk_clk),                                                                                      //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                                             // clk_reset.reset
		.in_data           (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                                          // (terminated)
		.csr_read          (1'b0),                                                                                                           // (terminated)
		.csr_write         (1'b0),                                                                                                           // (terminated)
		.csr_readdata      (),                                                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                           // (terminated)
		.almost_full_data  (),                                                                                                               // (terminated)
		.almost_empty_data (),                                                                                                               // (terminated)
		.in_startofpacket  (1'b0),                                                                                                           // (terminated)
		.in_endofpacket    (1'b0),                                                                                                           // (terminated)
		.out_startofpacket (),                                                                                                               // (terminated)
		.out_endofpacket   (),                                                                                                               // (terminated)
		.in_empty          (1'b0),                                                                                                           // (terminated)
		.out_empty         (),                                                                                                               // (terminated)
		.in_error          (1'b0),                                                                                                           // (terminated)
		.out_error         (),                                                                                                               // (terminated)
		.in_channel        (1'b0),                                                                                                           // (terminated)
		.out_channel       ()                                                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (80),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (87),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (95),
		.PKT_PROTECTION_L          (93),
		.PKT_RESPONSE_STATUS_H     (101),
		.PKT_RESPONSE_STATUS_L     (100),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.ST_CHANNEL_W              (20),
		.ST_DATA_W                 (102),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) i2c_scl_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c1_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src15_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src15_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src15_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src15_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src15_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src15_channel),                                                //                .channel
		.rf_sink_ready           (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (103),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c1_clk),                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (80),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (87),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (95),
		.PKT_PROTECTION_L          (93),
		.PKT_RESPONSE_STATUS_H     (101),
		.PKT_RESPONSE_STATUS_L     (100),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.ST_CHANNEL_W              (20),
		.ST_DATA_W                 (102),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) i2c_sda_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c1_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src16_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src16_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src16_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src16_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src16_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src16_channel),                                                //                .channel
		.rf_sink_ready           (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (103),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c1_clk),                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (80),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (87),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (95),
		.PKT_PROTECTION_L          (93),
		.PKT_RESPONSE_STATUS_H     (101),
		.PKT_RESPONSE_STATUS_L     (100),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.ST_CHANNEL_W              (20),
		.ST_DATA_W                 (102),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) i2c_scl_2_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c1_clk),                                                                   //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src17_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src17_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src17_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src17_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src17_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src17_channel),                                                  //                .channel
		.rf_sink_ready           (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (103),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c1_clk),                                                                   //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (80),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (87),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (95),
		.PKT_PROTECTION_L          (93),
		.PKT_RESPONSE_STATUS_H     (101),
		.PKT_RESPONSE_STATUS_L     (100),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.ST_CHANNEL_W              (20),
		.ST_DATA_W                 (102),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) i2c_sda_2_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c1_clk),                                                                   //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src18_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src18_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src18_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src18_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src18_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src18_channel),                                                  //                .channel
		.rf_sink_ready           (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (103),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c1_clk),                                                                   //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (80),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (87),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (95),
		.PKT_PROTECTION_L          (93),
		.PKT_RESPONSE_STATUS_H     (101),
		.PKT_RESPONSE_STATUS_L     (100),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.ST_CHANNEL_W              (20),
		.ST_DATA_W                 (102),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) drum_out_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c1_clk),                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                   //       clk_reset.reset
		.m0_address              (drum_out_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (drum_out_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (drum_out_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (drum_out_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (drum_out_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (drum_out_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (drum_out_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (drum_out_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (drum_out_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (drum_out_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (drum_out_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (drum_out_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (drum_out_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (drum_out_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (drum_out_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (drum_out_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src19_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src19_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src19_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src19_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src19_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src19_channel),                                                 //                .channel
		.rf_sink_ready           (drum_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (drum_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (drum_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (drum_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (drum_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (drum_out_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (drum_out_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (drum_out_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (drum_out_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (drum_out_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (drum_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (drum_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (drum_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (drum_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (drum_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (drum_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (103),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) drum_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c1_clk),                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.in_data           (drum_out_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (drum_out_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (drum_out_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (drum_out_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (drum_out_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (drum_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (drum_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (drum_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (drum_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (drum_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	niosII_system_addr_router addr_router (
		.sink_ready         (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                                             //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                       //       src.ready
		.src_valid          (addr_router_src_valid),                                                                       //          .valid
		.src_data           (addr_router_src_data),                                                                        //          .data
		.src_channel        (addr_router_src_channel),                                                                     //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                               //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                                  //          .endofpacket
	);

	niosII_system_addr_router_001 addr_router_001 (
		.sink_ready         (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                            //          .valid
		.src_data           (addr_router_001_src_data),                                                             //          .data
		.src_channel        (addr_router_001_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                       //          .endofpacket
	);

	niosII_system_id_router id_router (
		.sink_ready         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                       //       src.ready
		.src_valid          (id_router_src_valid),                                                                       //          .valid
		.src_data           (id_router_src_data),                                                                        //          .data
		.src_channel        (id_router_src_channel),                                                                     //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                               //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                                  //          .endofpacket
	);

	niosII_system_id_router id_router_001 (
		.sink_ready         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                        //       src.ready
		.src_valid          (id_router_001_src_valid),                                                        //          .valid
		.src_data           (id_router_001_src_data),                                                         //          .data
		.src_channel        (id_router_001_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                                   //          .endofpacket
	);

	niosII_system_id_router_002 id_router_002 (
		.sink_ready         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                               //       src.ready
		.src_valid          (id_router_002_src_valid),                                               //          .valid
		.src_data           (id_router_002_src_data),                                                //          .data
		.src_channel        (id_router_002_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                          //          .endofpacket
	);

	niosII_system_id_router_002 id_router_003 (
		.sink_ready         (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                      // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                             //       src.ready
		.src_valid          (id_router_003_src_valid),                                                             //          .valid
		.src_data           (id_router_003_src_data),                                                              //          .data
		.src_channel        (id_router_003_src_channel),                                                           //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                        //          .endofpacket
	);

	niosII_system_id_router id_router_004 (
		.sink_ready         (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sd_card_spi_master_spi_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                 // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                                        //       src.ready
		.src_valid          (id_router_004_src_valid),                                                                        //          .valid
		.src_data           (id_router_004_src_data),                                                                         //          .data
		.src_channel        (id_router_004_src_channel),                                                                      //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                                                //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                                   //          .endofpacket
	);

	niosII_system_id_router_005 id_router_005 (
		.sink_ready         (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (generic_tristate_controller_0_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                                      //       src.ready
		.src_valid          (id_router_005_src_valid),                                                                      //          .valid
		.src_data           (id_router_005_src_data),                                                                       //          .data
		.src_channel        (id_router_005_src_channel),                                                                    //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                                              //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                                                 //          .endofpacket
	);

	niosII_system_id_router_006 id_router_006 (
		.sink_ready         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                            // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                                       //       src.ready
		.src_valid          (id_router_006_src_valid),                                                       //          .valid
		.src_data           (id_router_006_src_data),                                                        //          .data
		.src_channel        (id_router_006_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                                  //          .endofpacket
	);

	niosII_system_id_router_006 id_router_007 (
		.sink_ready         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                                               //       src.ready
		.src_valid          (id_router_007_src_valid),                                                               //          .valid
		.src_data           (id_router_007_src_data),                                                                //          .data
		.src_channel        (id_router_007_src_channel),                                                             //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                                       //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                                          //          .endofpacket
	);

	niosII_system_id_router_006 id_router_008 (
		.sink_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                               //       src.ready
		.src_valid          (id_router_008_src_valid),                                               //          .valid
		.src_data           (id_router_008_src_data),                                                //          .data
		.src_channel        (id_router_008_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                          //          .endofpacket
	);

	niosII_system_id_router_006 id_router_009 (
		.sink_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_009_src_valid),                                                                  //          .valid
		.src_data           (id_router_009_src_data),                                                                   //          .data
		.src_channel        (id_router_009_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                                             //          .endofpacket
	);

	niosII_system_id_router_010 id_router_010 (
		.sink_ready         (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                                             //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                                                     //       src.ready
		.src_valid          (id_router_010_src_valid),                                                                     //          .valid
		.src_data           (id_router_010_src_data),                                                                      //          .data
		.src_channel        (id_router_010_src_channel),                                                                   //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                                             //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                                                //          .endofpacket
	);

	niosII_system_id_router_006 id_router_011 (
		.sink_ready         (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                                  //       src.ready
		.src_valid          (id_router_011_src_valid),                                                  //          .valid
		.src_data           (id_router_011_src_data),                                                   //          .data
		.src_channel        (id_router_011_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                             //          .endofpacket
	);

	niosII_system_id_router_006 id_router_012 (
		.sink_ready         (switch_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (switch_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (switch_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (switch_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (switch_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                                              //       src.ready
		.src_valid          (id_router_012_src_valid),                                              //          .valid
		.src_data           (id_router_012_src_data),                                               //          .data
		.src_channel        (id_router_012_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)                                         //          .endofpacket
	);

	niosII_system_id_router_006 id_router_013 (
		.sink_ready         (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (up_clocks_1_audio_clk_clk),                                                             //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (id_router_013_src_ready),                                                               //       src.ready
		.src_valid          (id_router_013_src_valid),                                                               //          .valid
		.src_data           (id_router_013_src_data),                                                                //          .data
		.src_channel        (id_router_013_src_channel),                                                             //          .channel
		.src_startofpacket  (id_router_013_src_startofpacket),                                                       //          .startofpacket
		.src_endofpacket    (id_router_013_src_endofpacket)                                                          //          .endofpacket
	);

	niosII_system_id_router_006 id_router_014 (
		.sink_ready         (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (up_clocks_1_audio_clk_clk),                                                                                  //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                                                         // clk_reset.reset
		.src_ready          (id_router_014_src_ready),                                                                                    //       src.ready
		.src_valid          (id_router_014_src_valid),                                                                                    //          .valid
		.src_data           (id_router_014_src_data),                                                                                     //          .data
		.src_channel        (id_router_014_src_channel),                                                                                  //          .channel
		.src_startofpacket  (id_router_014_src_startofpacket),                                                                            //          .startofpacket
		.src_endofpacket    (id_router_014_src_endofpacket)                                                                               //          .endofpacket
	);

	niosII_system_id_router_006 id_router_015 (
		.sink_ready         (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_015_src_ready),                                               //       src.ready
		.src_valid          (id_router_015_src_valid),                                               //          .valid
		.src_data           (id_router_015_src_data),                                                //          .data
		.src_channel        (id_router_015_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_015_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_015_src_endofpacket)                                          //          .endofpacket
	);

	niosII_system_id_router_006 id_router_016 (
		.sink_ready         (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_016_src_ready),                                               //       src.ready
		.src_valid          (id_router_016_src_valid),                                               //          .valid
		.src_data           (id_router_016_src_data),                                                //          .data
		.src_channel        (id_router_016_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_016_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_016_src_endofpacket)                                          //          .endofpacket
	);

	niosII_system_id_router_006 id_router_017 (
		.sink_ready         (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (i2c_scl_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_017_src_ready),                                                 //       src.ready
		.src_valid          (id_router_017_src_valid),                                                 //          .valid
		.src_data           (id_router_017_src_data),                                                  //          .data
		.src_channel        (id_router_017_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_017_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_017_src_endofpacket)                                            //          .endofpacket
	);

	niosII_system_id_router_006 id_router_018 (
		.sink_ready         (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (i2c_sda_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_018_src_ready),                                                 //       src.ready
		.src_valid          (id_router_018_src_valid),                                                 //          .valid
		.src_data           (id_router_018_src_data),                                                  //          .data
		.src_channel        (id_router_018_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_018_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_018_src_endofpacket)                                            //          .endofpacket
	);

	niosII_system_id_router_006 id_router_019 (
		.sink_ready         (drum_out_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (drum_out_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (drum_out_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (drum_out_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (drum_out_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                         // clk_reset.reset
		.src_ready          (id_router_019_src_ready),                                                //       src.ready
		.src_valid          (id_router_019_src_valid),                                                //          .valid
		.src_data           (id_router_019_src_data),                                                 //          .data
		.src_channel        (id_router_019_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_019_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_019_src_endofpacket)                                           //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (87),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.MAX_OUTSTANDING_RESPONSES (9),
		.PIPELINED                 (0),
		.ST_DATA_W                 (102),
		.ST_CHANNEL_W              (20),
		.VALID_WIDTH               (20),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (altpll_0_c1_clk),                //       clk.clk
		.reset                  (rst_controller_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_src_data),           //          .data
		.cmd_sink_channel       (addr_router_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (87),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.MAX_OUTSTANDING_RESPONSES (9),
		.PIPELINED                 (0),
		.ST_DATA_W                 (102),
		.ST_CHANNEL_W              (20),
		.VALID_WIDTH               (20),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_001 (
		.clk                    (altpll_0_c1_clk),                    //       clk.clk
		.reset                  (rst_controller_reset_out_reset),     // clk_reset.reset
		.cmd_sink_ready         (addr_router_001_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_001_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_001_src_data),           //          .data
		.cmd_sink_channel       (addr_router_001_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_001_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_001_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_001_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_001_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_001_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_001_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_001_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_001_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_001_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_001_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_001_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_001_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_001_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_001_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_001_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_001_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_001_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_001_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_001_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_001_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (42),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (62),
		.PKT_BYTE_CNT_H            (51),
		.PKT_BYTE_CNT_L            (49),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (57),
		.PKT_BURST_SIZE_L          (55),
		.PKT_BURST_TYPE_H          (59),
		.PKT_BURST_TYPE_L          (58),
		.PKT_BURSTWRAP_H           (54),
		.PKT_BURSTWRAP_L           (52),
		.PKT_TRANS_COMPRESSED_READ (43),
		.PKT_TRANS_WRITE           (45),
		.PKT_TRANS_READ            (46),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (84),
		.ST_CHANNEL_W              (20),
		.OUT_BYTE_CNT_H            (50),
		.OUT_BURSTWRAP_H           (54),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter (
		.clk                   (altpll_0_c1_clk),                     //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (width_adapter_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_src_data),              //          .data
		.sink0_channel         (width_adapter_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_src_ready),             //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (42),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (62),
		.PKT_BYTE_CNT_H            (51),
		.PKT_BYTE_CNT_L            (49),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (57),
		.PKT_BURST_SIZE_L          (55),
		.PKT_BURST_TYPE_H          (59),
		.PKT_BURST_TYPE_L          (58),
		.PKT_BURSTWRAP_H           (54),
		.PKT_BURSTWRAP_L           (52),
		.PKT_TRANS_COMPRESSED_READ (43),
		.PKT_TRANS_WRITE           (45),
		.PKT_TRANS_READ            (46),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (84),
		.ST_CHANNEL_W              (20),
		.OUT_BYTE_CNT_H            (50),
		.OUT_BURSTWRAP_H           (54),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter_001 (
		.clk                   (altpll_0_c1_clk),                         //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (width_adapter_002_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_002_src_data),              //          .data
		.sink0_channel         (width_adapter_002_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_002_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_002_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_002_src_ready),             //          .ready
		.source0_valid         (burst_adapter_001_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_001_source0_data),          //          .data
		.source0_channel       (burst_adapter_001_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_001_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_001_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_001_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (33),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (53),
		.PKT_BYTE_CNT_H            (42),
		.PKT_BYTE_CNT_L            (40),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURST_SIZE_H          (48),
		.PKT_BURST_SIZE_L          (46),
		.PKT_BURST_TYPE_H          (50),
		.PKT_BURST_TYPE_L          (49),
		.PKT_BURSTWRAP_H           (45),
		.PKT_BURSTWRAP_L           (43),
		.PKT_TRANS_COMPRESSED_READ (34),
		.PKT_TRANS_WRITE           (36),
		.PKT_TRANS_READ            (37),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (75),
		.ST_CHANNEL_W              (20),
		.OUT_BYTE_CNT_H            (40),
		.OUT_BURSTWRAP_H           (45),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter_002 (
		.clk                   (altpll_0_c1_clk),                         //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (width_adapter_004_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_004_src_data),              //          .data
		.sink0_channel         (width_adapter_004_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_004_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_004_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_004_src_ready),             //          .ready
		.source0_valid         (burst_adapter_002_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_002_source0_data),          //          .data
		.source0_channel       (burst_adapter_002_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_002_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_002_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_002_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (33),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (53),
		.PKT_BYTE_CNT_H            (42),
		.PKT_BYTE_CNT_L            (40),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURST_SIZE_H          (48),
		.PKT_BURST_SIZE_L          (46),
		.PKT_BURST_TYPE_H          (50),
		.PKT_BURST_TYPE_L          (49),
		.PKT_BURSTWRAP_H           (45),
		.PKT_BURSTWRAP_L           (43),
		.PKT_TRANS_COMPRESSED_READ (34),
		.PKT_TRANS_WRITE           (36),
		.PKT_TRANS_READ            (37),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (75),
		.ST_CHANNEL_W              (20),
		.OUT_BYTE_CNT_H            (40),
		.OUT_BURSTWRAP_H           (45),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_003 (
		.clk                   (altpll_0_c1_clk),                         //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (width_adapter_006_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_006_src_data),              //          .data
		.sink0_channel         (width_adapter_006_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_006_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_006_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_006_src_ready),             //          .ready
		.source0_valid         (burst_adapter_003_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_003_source0_data),          //          .data
		.source0_channel       (burst_adapter_003_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_003_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_003_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_003_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in0.reset
		.reset_in1  (~reset_reset_n),                             // reset_in1.reset
		.clk        (altpll_0_c1_clk),                            //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),             // reset_out.reset
		.reset_in2  (1'b0),                                       // (terminated)
		.reset_in3  (1'b0),                                       // (terminated)
		.reset_in4  (1'b0),                                       // (terminated)
		.reset_in5  (1'b0),                                       // (terminated)
		.reset_in6  (1'b0),                                       // (terminated)
		.reset_in7  (1'b0),                                       // (terminated)
		.reset_in8  (1'b0),                                       // (terminated)
		.reset_in9  (1'b0),                                       // (terminated)
		.reset_in10 (1'b0),                                       // (terminated)
		.reset_in11 (1'b0),                                       // (terminated)
		.reset_in12 (1'b0),                                       // (terminated)
		.reset_in13 (1'b0),                                       // (terminated)
		.reset_in14 (1'b0),                                       // (terminated)
		.reset_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_001 (
		.reset_in0  (~reset_reset_n),                             // reset_in0.reset
		.reset_in1  (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clk_clk),                                    //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset),         // reset_out.reset
		.reset_in2  (1'b0),                                       // (terminated)
		.reset_in3  (1'b0),                                       // (terminated)
		.reset_in4  (1'b0),                                       // (terminated)
		.reset_in5  (1'b0),                                       // (terminated)
		.reset_in6  (1'b0),                                       // (terminated)
		.reset_in7  (1'b0),                                       // (terminated)
		.reset_in8  (1'b0),                                       // (terminated)
		.reset_in9  (1'b0),                                       // (terminated)
		.reset_in10 (1'b0),                                       // (terminated)
		.reset_in11 (1'b0),                                       // (terminated)
		.reset_in12 (1'b0),                                       // (terminated)
		.reset_in13 (1'b0),                                       // (terminated)
		.reset_in14 (1'b0),                                       // (terminated)
		.reset_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_002 (
		.reset_in0  (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in0.reset
		.reset_in1  (~reset_reset_n),                             // reset_in1.reset
		.clk        (up_clocks_1_audio_clk_clk),                  //       clk.clk
		.reset_out  (rst_controller_002_reset_out_reset),         // reset_out.reset
		.reset_in2  (1'b0),                                       // (terminated)
		.reset_in3  (1'b0),                                       // (terminated)
		.reset_in4  (1'b0),                                       // (terminated)
		.reset_in5  (1'b0),                                       // (terminated)
		.reset_in6  (1'b0),                                       // (terminated)
		.reset_in7  (1'b0),                                       // (terminated)
		.reset_in8  (1'b0),                                       // (terminated)
		.reset_in9  (1'b0),                                       // (terminated)
		.reset_in10 (1'b0),                                       // (terminated)
		.reset_in11 (1'b0),                                       // (terminated)
		.reset_in12 (1'b0),                                       // (terminated)
		.reset_in13 (1'b0),                                       // (terminated)
		.reset_in14 (1'b0),                                       // (terminated)
		.reset_in15 (1'b0)                                        // (terminated)
	);

	niosII_system_cmd_xbar_demux cmd_xbar_demux (
		.clk                (altpll_0_c1_clk),                   //        clk.clk
		.reset              (rst_controller_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),           //           .channel
		.sink_data          (limiter_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket),   //           .endofpacket
		.src3_ready         (cmd_xbar_demux_src3_ready),         //       src3.ready
		.src3_valid         (cmd_xbar_demux_src3_valid),         //           .valid
		.src3_data          (cmd_xbar_demux_src3_data),          //           .data
		.src3_channel       (cmd_xbar_demux_src3_channel),       //           .channel
		.src3_startofpacket (cmd_xbar_demux_src3_startofpacket), //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_src3_endofpacket),   //           .endofpacket
		.src4_ready         (cmd_xbar_demux_src4_ready),         //       src4.ready
		.src4_valid         (cmd_xbar_demux_src4_valid),         //           .valid
		.src4_data          (cmd_xbar_demux_src4_data),          //           .data
		.src4_channel       (cmd_xbar_demux_src4_channel),       //           .channel
		.src4_startofpacket (cmd_xbar_demux_src4_startofpacket), //           .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_src4_endofpacket),   //           .endofpacket
		.src5_ready         (cmd_xbar_demux_src5_ready),         //       src5.ready
		.src5_valid         (cmd_xbar_demux_src5_valid),         //           .valid
		.src5_data          (cmd_xbar_demux_src5_data),          //           .data
		.src5_channel       (cmd_xbar_demux_src5_channel),       //           .channel
		.src5_startofpacket (cmd_xbar_demux_src5_startofpacket), //           .startofpacket
		.src5_endofpacket   (cmd_xbar_demux_src5_endofpacket)    //           .endofpacket
	);

	niosII_system_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                 (altpll_0_c1_clk),                        //        clk.clk
		.reset               (rst_controller_reset_out_reset),         //  clk_reset.reset
		.sink_ready          (limiter_001_cmd_src_ready),              //       sink.ready
		.sink_channel        (limiter_001_cmd_src_channel),            //           .channel
		.sink_data           (limiter_001_cmd_src_data),               //           .data
		.sink_startofpacket  (limiter_001_cmd_src_startofpacket),      //           .startofpacket
		.sink_endofpacket    (limiter_001_cmd_src_endofpacket),        //           .endofpacket
		.sink_valid          (limiter_001_cmd_valid_data),             // sink_valid.data
		.src0_ready          (cmd_xbar_demux_001_src0_ready),          //       src0.ready
		.src0_valid          (cmd_xbar_demux_001_src0_valid),          //           .valid
		.src0_data           (cmd_xbar_demux_001_src0_data),           //           .data
		.src0_channel        (cmd_xbar_demux_001_src0_channel),        //           .channel
		.src0_startofpacket  (cmd_xbar_demux_001_src0_startofpacket),  //           .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_001_src0_endofpacket),    //           .endofpacket
		.src1_ready          (cmd_xbar_demux_001_src1_ready),          //       src1.ready
		.src1_valid          (cmd_xbar_demux_001_src1_valid),          //           .valid
		.src1_data           (cmd_xbar_demux_001_src1_data),           //           .data
		.src1_channel        (cmd_xbar_demux_001_src1_channel),        //           .channel
		.src1_startofpacket  (cmd_xbar_demux_001_src1_startofpacket),  //           .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_001_src1_endofpacket),    //           .endofpacket
		.src2_ready          (cmd_xbar_demux_001_src2_ready),          //       src2.ready
		.src2_valid          (cmd_xbar_demux_001_src2_valid),          //           .valid
		.src2_data           (cmd_xbar_demux_001_src2_data),           //           .data
		.src2_channel        (cmd_xbar_demux_001_src2_channel),        //           .channel
		.src2_startofpacket  (cmd_xbar_demux_001_src2_startofpacket),  //           .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_001_src2_endofpacket),    //           .endofpacket
		.src3_ready          (cmd_xbar_demux_001_src3_ready),          //       src3.ready
		.src3_valid          (cmd_xbar_demux_001_src3_valid),          //           .valid
		.src3_data           (cmd_xbar_demux_001_src3_data),           //           .data
		.src3_channel        (cmd_xbar_demux_001_src3_channel),        //           .channel
		.src3_startofpacket  (cmd_xbar_demux_001_src3_startofpacket),  //           .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_001_src3_endofpacket),    //           .endofpacket
		.src4_ready          (cmd_xbar_demux_001_src4_ready),          //       src4.ready
		.src4_valid          (cmd_xbar_demux_001_src4_valid),          //           .valid
		.src4_data           (cmd_xbar_demux_001_src4_data),           //           .data
		.src4_channel        (cmd_xbar_demux_001_src4_channel),        //           .channel
		.src4_startofpacket  (cmd_xbar_demux_001_src4_startofpacket),  //           .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_001_src4_endofpacket),    //           .endofpacket
		.src5_ready          (cmd_xbar_demux_001_src5_ready),          //       src5.ready
		.src5_valid          (cmd_xbar_demux_001_src5_valid),          //           .valid
		.src5_data           (cmd_xbar_demux_001_src5_data),           //           .data
		.src5_channel        (cmd_xbar_demux_001_src5_channel),        //           .channel
		.src5_startofpacket  (cmd_xbar_demux_001_src5_startofpacket),  //           .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_001_src5_endofpacket),    //           .endofpacket
		.src6_ready          (cmd_xbar_demux_001_src6_ready),          //       src6.ready
		.src6_valid          (cmd_xbar_demux_001_src6_valid),          //           .valid
		.src6_data           (cmd_xbar_demux_001_src6_data),           //           .data
		.src6_channel        (cmd_xbar_demux_001_src6_channel),        //           .channel
		.src6_startofpacket  (cmd_xbar_demux_001_src6_startofpacket),  //           .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_001_src6_endofpacket),    //           .endofpacket
		.src7_ready          (cmd_xbar_demux_001_src7_ready),          //       src7.ready
		.src7_valid          (cmd_xbar_demux_001_src7_valid),          //           .valid
		.src7_data           (cmd_xbar_demux_001_src7_data),           //           .data
		.src7_channel        (cmd_xbar_demux_001_src7_channel),        //           .channel
		.src7_startofpacket  (cmd_xbar_demux_001_src7_startofpacket),  //           .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_001_src7_endofpacket),    //           .endofpacket
		.src8_ready          (cmd_xbar_demux_001_src8_ready),          //       src8.ready
		.src8_valid          (cmd_xbar_demux_001_src8_valid),          //           .valid
		.src8_data           (cmd_xbar_demux_001_src8_data),           //           .data
		.src8_channel        (cmd_xbar_demux_001_src8_channel),        //           .channel
		.src8_startofpacket  (cmd_xbar_demux_001_src8_startofpacket),  //           .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_001_src8_endofpacket),    //           .endofpacket
		.src9_ready          (cmd_xbar_demux_001_src9_ready),          //       src9.ready
		.src9_valid          (cmd_xbar_demux_001_src9_valid),          //           .valid
		.src9_data           (cmd_xbar_demux_001_src9_data),           //           .data
		.src9_channel        (cmd_xbar_demux_001_src9_channel),        //           .channel
		.src9_startofpacket  (cmd_xbar_demux_001_src9_startofpacket),  //           .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_001_src9_endofpacket),    //           .endofpacket
		.src10_ready         (cmd_xbar_demux_001_src10_ready),         //      src10.ready
		.src10_valid         (cmd_xbar_demux_001_src10_valid),         //           .valid
		.src10_data          (cmd_xbar_demux_001_src10_data),          //           .data
		.src10_channel       (cmd_xbar_demux_001_src10_channel),       //           .channel
		.src10_startofpacket (cmd_xbar_demux_001_src10_startofpacket), //           .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_001_src10_endofpacket),   //           .endofpacket
		.src11_ready         (cmd_xbar_demux_001_src11_ready),         //      src11.ready
		.src11_valid         (cmd_xbar_demux_001_src11_valid),         //           .valid
		.src11_data          (cmd_xbar_demux_001_src11_data),          //           .data
		.src11_channel       (cmd_xbar_demux_001_src11_channel),       //           .channel
		.src11_startofpacket (cmd_xbar_demux_001_src11_startofpacket), //           .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_001_src11_endofpacket),   //           .endofpacket
		.src12_ready         (cmd_xbar_demux_001_src12_ready),         //      src12.ready
		.src12_valid         (cmd_xbar_demux_001_src12_valid),         //           .valid
		.src12_data          (cmd_xbar_demux_001_src12_data),          //           .data
		.src12_channel       (cmd_xbar_demux_001_src12_channel),       //           .channel
		.src12_startofpacket (cmd_xbar_demux_001_src12_startofpacket), //           .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_001_src12_endofpacket),   //           .endofpacket
		.src13_ready         (cmd_xbar_demux_001_src13_ready),         //      src13.ready
		.src13_valid         (cmd_xbar_demux_001_src13_valid),         //           .valid
		.src13_data          (cmd_xbar_demux_001_src13_data),          //           .data
		.src13_channel       (cmd_xbar_demux_001_src13_channel),       //           .channel
		.src13_startofpacket (cmd_xbar_demux_001_src13_startofpacket), //           .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_001_src13_endofpacket),   //           .endofpacket
		.src14_ready         (cmd_xbar_demux_001_src14_ready),         //      src14.ready
		.src14_valid         (cmd_xbar_demux_001_src14_valid),         //           .valid
		.src14_data          (cmd_xbar_demux_001_src14_data),          //           .data
		.src14_channel       (cmd_xbar_demux_001_src14_channel),       //           .channel
		.src14_startofpacket (cmd_xbar_demux_001_src14_startofpacket), //           .startofpacket
		.src14_endofpacket   (cmd_xbar_demux_001_src14_endofpacket),   //           .endofpacket
		.src15_ready         (cmd_xbar_demux_001_src15_ready),         //      src15.ready
		.src15_valid         (cmd_xbar_demux_001_src15_valid),         //           .valid
		.src15_data          (cmd_xbar_demux_001_src15_data),          //           .data
		.src15_channel       (cmd_xbar_demux_001_src15_channel),       //           .channel
		.src15_startofpacket (cmd_xbar_demux_001_src15_startofpacket), //           .startofpacket
		.src15_endofpacket   (cmd_xbar_demux_001_src15_endofpacket),   //           .endofpacket
		.src16_ready         (cmd_xbar_demux_001_src16_ready),         //      src16.ready
		.src16_valid         (cmd_xbar_demux_001_src16_valid),         //           .valid
		.src16_data          (cmd_xbar_demux_001_src16_data),          //           .data
		.src16_channel       (cmd_xbar_demux_001_src16_channel),       //           .channel
		.src16_startofpacket (cmd_xbar_demux_001_src16_startofpacket), //           .startofpacket
		.src16_endofpacket   (cmd_xbar_demux_001_src16_endofpacket),   //           .endofpacket
		.src17_ready         (cmd_xbar_demux_001_src17_ready),         //      src17.ready
		.src17_valid         (cmd_xbar_demux_001_src17_valid),         //           .valid
		.src17_data          (cmd_xbar_demux_001_src17_data),          //           .data
		.src17_channel       (cmd_xbar_demux_001_src17_channel),       //           .channel
		.src17_startofpacket (cmd_xbar_demux_001_src17_startofpacket), //           .startofpacket
		.src17_endofpacket   (cmd_xbar_demux_001_src17_endofpacket),   //           .endofpacket
		.src18_ready         (cmd_xbar_demux_001_src18_ready),         //      src18.ready
		.src18_valid         (cmd_xbar_demux_001_src18_valid),         //           .valid
		.src18_data          (cmd_xbar_demux_001_src18_data),          //           .data
		.src18_channel       (cmd_xbar_demux_001_src18_channel),       //           .channel
		.src18_startofpacket (cmd_xbar_demux_001_src18_startofpacket), //           .startofpacket
		.src18_endofpacket   (cmd_xbar_demux_001_src18_endofpacket),   //           .endofpacket
		.src19_ready         (cmd_xbar_demux_001_src19_ready),         //      src19.ready
		.src19_valid         (cmd_xbar_demux_001_src19_valid),         //           .valid
		.src19_data          (cmd_xbar_demux_001_src19_data),          //           .data
		.src19_channel       (cmd_xbar_demux_001_src19_channel),       //           .channel
		.src19_startofpacket (cmd_xbar_demux_001_src19_startofpacket), //           .startofpacket
		.src19_endofpacket   (cmd_xbar_demux_001_src19_endofpacket)    //           .endofpacket
	);

	niosII_system_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (altpll_0_c1_clk),                       //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (altpll_0_c1_clk),                       //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	niosII_system_cmd_xbar_mux cmd_xbar_mux_002 (
		.clk                 (altpll_0_c1_clk),                       //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src2_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src2_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src2_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src2_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src2_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src2_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src2_endofpacket)    //          .endofpacket
	);

	niosII_system_cmd_xbar_mux cmd_xbar_mux_003 (
		.clk                 (altpll_0_c1_clk),                       //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_003_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_003_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_003_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_003_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_003_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_003_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src3_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src3_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src3_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src3_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src3_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src3_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src3_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src3_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src3_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src3_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src3_endofpacket)    //          .endofpacket
	);

	niosII_system_cmd_xbar_mux cmd_xbar_mux_004 (
		.clk                 (altpll_0_c1_clk),                       //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_004_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_004_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_004_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_004_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_004_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_004_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src4_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src4_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src4_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src4_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src4_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src4_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src4_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src4_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src4_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src4_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src4_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src4_endofpacket)    //          .endofpacket
	);

	niosII_system_cmd_xbar_mux cmd_xbar_mux_005 (
		.clk                 (altpll_0_c1_clk),                       //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_005_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_005_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_005_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_005_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_005_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_005_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src5_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src5_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src5_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src5_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src5_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src5_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src5_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src5_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src5_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src5_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src5_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src5_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux rsp_xbar_demux (
		.clk                (altpll_0_c1_clk),                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (altpll_0_c1_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux rsp_xbar_demux_002 (
		.clk                (altpll_0_c1_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (width_adapter_001_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_001_src_channel),         //          .channel
		.sink_data          (width_adapter_001_src_data),            //          .data
		.sink_startofpacket (width_adapter_001_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_001_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_001_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux rsp_xbar_demux_003 (
		.clk                (altpll_0_c1_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (width_adapter_003_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_003_src_channel),         //          .channel
		.sink_data          (width_adapter_003_src_data),            //          .data
		.sink_startofpacket (width_adapter_003_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_003_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_003_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_003_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_003_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_003_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_003_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_003_src1_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux rsp_xbar_demux_004 (
		.clk                (altpll_0_c1_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_004_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_004_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_004_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_004_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_004_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_004_src1_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux rsp_xbar_demux_005 (
		.clk                (altpll_0_c1_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (width_adapter_005_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_005_src_channel),         //          .channel
		.sink_data          (width_adapter_005_src_data),            //          .data
		.sink_startofpacket (width_adapter_005_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_005_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_005_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_005_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_005_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_005_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_005_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_005_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_005_src1_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_006 rsp_xbar_demux_006 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_006 rsp_xbar_demux_007 (
		.clk                (altpll_0_c1_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_006 rsp_xbar_demux_008 (
		.clk                (altpll_0_c1_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_006 rsp_xbar_demux_009 (
		.clk                (altpll_0_c1_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_006 rsp_xbar_demux_010 (
		.clk                (altpll_0_c1_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (width_adapter_007_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_007_src_channel),         //          .channel
		.sink_data          (width_adapter_007_src_data),            //          .data
		.sink_startofpacket (width_adapter_007_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_007_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_007_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_006 rsp_xbar_demux_011 (
		.clk                (altpll_0_c1_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_011_src_ready),               //      sink.ready
		.sink_channel       (id_router_011_src_channel),             //          .channel
		.sink_data          (id_router_011_src_data),                //          .data
		.sink_startofpacket (id_router_011_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_011_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_011_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_006 rsp_xbar_demux_012 (
		.clk                (altpll_0_c1_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_012_src_ready),               //      sink.ready
		.sink_channel       (id_router_012_src_channel),             //          .channel
		.sink_data          (id_router_012_src_data),                //          .data
		.sink_startofpacket (id_router_012_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_012_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_012_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_006 rsp_xbar_demux_013 (
		.clk                (up_clocks_1_audio_clk_clk),             //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_013_src_ready),               //      sink.ready
		.sink_channel       (id_router_013_src_channel),             //          .channel
		.sink_data          (id_router_013_src_data),                //          .data
		.sink_startofpacket (id_router_013_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_013_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_013_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_013_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_013_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_006 rsp_xbar_demux_014 (
		.clk                (up_clocks_1_audio_clk_clk),             //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_014_src_ready),               //      sink.ready
		.sink_channel       (id_router_014_src_channel),             //          .channel
		.sink_data          (id_router_014_src_data),                //          .data
		.sink_startofpacket (id_router_014_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_014_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_014_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_014_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_014_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_006 rsp_xbar_demux_015 (
		.clk                (altpll_0_c1_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_015_src_ready),               //      sink.ready
		.sink_channel       (id_router_015_src_channel),             //          .channel
		.sink_data          (id_router_015_src_data),                //          .data
		.sink_startofpacket (id_router_015_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_015_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_015_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_015_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_015_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_006 rsp_xbar_demux_016 (
		.clk                (altpll_0_c1_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_016_src_ready),               //      sink.ready
		.sink_channel       (id_router_016_src_channel),             //          .channel
		.sink_data          (id_router_016_src_data),                //          .data
		.sink_startofpacket (id_router_016_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_016_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_016_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_016_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_016_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_006 rsp_xbar_demux_017 (
		.clk                (altpll_0_c1_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_017_src_ready),               //      sink.ready
		.sink_channel       (id_router_017_src_channel),             //          .channel
		.sink_data          (id_router_017_src_data),                //          .data
		.sink_startofpacket (id_router_017_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_017_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_017_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_017_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_017_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_006 rsp_xbar_demux_018 (
		.clk                (altpll_0_c1_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_018_src_ready),               //      sink.ready
		.sink_channel       (id_router_018_src_channel),             //          .channel
		.sink_data          (id_router_018_src_data),                //          .data
		.sink_startofpacket (id_router_018_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_018_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_018_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_018_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_018_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_006 rsp_xbar_demux_019 (
		.clk                (altpll_0_c1_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_019_src_ready),               //      sink.ready
		.sink_channel       (id_router_019_src_channel),             //          .channel
		.sink_data          (id_router_019_src_data),                //          .data
		.sink_startofpacket (id_router_019_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_019_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_019_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_019_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_019_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_019_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_019_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_019_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (altpll_0_c1_clk),                       //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready         (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                  (altpll_0_c1_clk),                       //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready            (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel        (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data           (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket  (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_002_src1_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_002_src1_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_002_src1_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_002_src1_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_003_src1_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_003_src1_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_003_src1_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_003_src1_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_003_src1_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_004_src1_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_004_src1_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_004_src1_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_004_src1_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_004_src1_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_004_src1_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_005_src1_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_005_src1_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_005_src1_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_005_src1_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_005_src1_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_005_src1_endofpacket),   //          .endofpacket
		.sink6_ready          (crosser_003_out_ready),                 //     sink6.ready
		.sink6_valid          (crosser_003_out_valid),                 //          .valid
		.sink6_channel        (crosser_003_out_channel),               //          .channel
		.sink6_data           (crosser_003_out_data),                  //          .data
		.sink6_startofpacket  (crosser_003_out_startofpacket),         //          .startofpacket
		.sink6_endofpacket    (crosser_003_out_endofpacket),           //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_008_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_008_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_009_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_009_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_010_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_011_src0_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_011_src0_endofpacket),   //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_012_src0_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_012_src0_endofpacket),   //          .endofpacket
		.sink13_ready         (crosser_004_out_ready),                 //    sink13.ready
		.sink13_valid         (crosser_004_out_valid),                 //          .valid
		.sink13_channel       (crosser_004_out_channel),               //          .channel
		.sink13_data          (crosser_004_out_data),                  //          .data
		.sink13_startofpacket (crosser_004_out_startofpacket),         //          .startofpacket
		.sink13_endofpacket   (crosser_004_out_endofpacket),           //          .endofpacket
		.sink14_ready         (crosser_005_out_ready),                 //    sink14.ready
		.sink14_valid         (crosser_005_out_valid),                 //          .valid
		.sink14_channel       (crosser_005_out_channel),               //          .channel
		.sink14_data          (crosser_005_out_data),                  //          .data
		.sink14_startofpacket (crosser_005_out_startofpacket),         //          .startofpacket
		.sink14_endofpacket   (crosser_005_out_endofpacket),           //          .endofpacket
		.sink15_ready         (rsp_xbar_demux_015_src0_ready),         //    sink15.ready
		.sink15_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.sink15_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.sink15_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.sink15_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.sink15_endofpacket   (rsp_xbar_demux_015_src0_endofpacket),   //          .endofpacket
		.sink16_ready         (rsp_xbar_demux_016_src0_ready),         //    sink16.ready
		.sink16_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.sink16_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.sink16_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.sink16_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.sink16_endofpacket   (rsp_xbar_demux_016_src0_endofpacket),   //          .endofpacket
		.sink17_ready         (rsp_xbar_demux_017_src0_ready),         //    sink17.ready
		.sink17_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.sink17_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.sink17_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.sink17_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.sink17_endofpacket   (rsp_xbar_demux_017_src0_endofpacket),   //          .endofpacket
		.sink18_ready         (rsp_xbar_demux_018_src0_ready),         //    sink18.ready
		.sink18_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.sink18_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.sink18_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.sink18_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.sink18_endofpacket   (rsp_xbar_demux_018_src0_endofpacket),   //          .endofpacket
		.sink19_ready         (rsp_xbar_demux_019_src0_ready),         //    sink19.ready
		.sink19_valid         (rsp_xbar_demux_019_src0_valid),         //          .valid
		.sink19_channel       (rsp_xbar_demux_019_src0_channel),       //          .channel
		.sink19_data          (rsp_xbar_demux_019_src0_data),          //          .data
		.sink19_startofpacket (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.sink19_endofpacket   (rsp_xbar_demux_019_src0_endofpacket)    //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (60),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (69),
		.IN_PKT_BYTE_CNT_L             (67),
		.IN_PKT_TRANS_COMPRESSED_READ  (61),
		.IN_PKT_BURSTWRAP_H            (72),
		.IN_PKT_BURSTWRAP_L            (70),
		.IN_PKT_BURST_SIZE_H           (75),
		.IN_PKT_BURST_SIZE_L           (73),
		.IN_PKT_RESPONSE_STATUS_H      (101),
		.IN_PKT_RESPONSE_STATUS_L      (100),
		.IN_PKT_TRANS_EXCLUSIVE        (66),
		.IN_PKT_BURST_TYPE_H           (77),
		.IN_PKT_BURST_TYPE_L           (76),
		.IN_ST_DATA_W                  (102),
		.OUT_PKT_ADDR_H                (42),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (51),
		.OUT_PKT_BYTE_CNT_L            (49),
		.OUT_PKT_TRANS_COMPRESSED_READ (43),
		.OUT_PKT_BURST_SIZE_H          (57),
		.OUT_PKT_BURST_SIZE_L          (55),
		.OUT_PKT_RESPONSE_STATUS_H     (83),
		.OUT_PKT_RESPONSE_STATUS_L     (82),
		.OUT_PKT_TRANS_EXCLUSIVE       (48),
		.OUT_PKT_BURST_TYPE_H          (59),
		.OUT_PKT_BURST_TYPE_L          (58),
		.OUT_ST_DATA_W                 (84),
		.ST_CHANNEL_W                  (20),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter (
		.clk                  (altpll_0_c1_clk),                    //       clk.clk
		.reset                (rst_controller_reset_out_reset),     // clk_reset.reset
		.in_valid             (cmd_xbar_mux_002_src_valid),         //      sink.valid
		.in_channel           (cmd_xbar_mux_002_src_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_mux_002_src_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_mux_002_src_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_mux_002_src_ready),         //          .ready
		.in_data              (cmd_xbar_mux_002_src_data),          //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),      //       src.endofpacket
		.out_data             (width_adapter_src_data),             //          .data
		.out_channel          (width_adapter_src_channel),          //          .channel
		.out_valid            (width_adapter_src_valid),            //          .valid
		.out_ready            (width_adapter_src_ready),            //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),    //          .startofpacket
		.in_command_size_data (3'b000)                              // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (42),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (51),
		.IN_PKT_BYTE_CNT_L             (49),
		.IN_PKT_TRANS_COMPRESSED_READ  (43),
		.IN_PKT_BURSTWRAP_H            (54),
		.IN_PKT_BURSTWRAP_L            (52),
		.IN_PKT_BURST_SIZE_H           (57),
		.IN_PKT_BURST_SIZE_L           (55),
		.IN_PKT_RESPONSE_STATUS_H      (83),
		.IN_PKT_RESPONSE_STATUS_L      (82),
		.IN_PKT_TRANS_EXCLUSIVE        (48),
		.IN_PKT_BURST_TYPE_H           (59),
		.IN_PKT_BURST_TYPE_L           (58),
		.IN_ST_DATA_W                  (84),
		.OUT_PKT_ADDR_H                (60),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (69),
		.OUT_PKT_BYTE_CNT_L            (67),
		.OUT_PKT_TRANS_COMPRESSED_READ (61),
		.OUT_PKT_BURST_SIZE_H          (75),
		.OUT_PKT_BURST_SIZE_L          (73),
		.OUT_PKT_RESPONSE_STATUS_H     (101),
		.OUT_PKT_RESPONSE_STATUS_L     (100),
		.OUT_PKT_TRANS_EXCLUSIVE       (66),
		.OUT_PKT_BURST_TYPE_H          (77),
		.OUT_PKT_BURST_TYPE_L          (76),
		.OUT_ST_DATA_W                 (102),
		.ST_CHANNEL_W                  (20),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_001 (
		.clk                  (altpll_0_c1_clk),                     //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (id_router_002_src_valid),             //      sink.valid
		.in_channel           (id_router_002_src_channel),           //          .channel
		.in_startofpacket     (id_router_002_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_002_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_002_src_ready),             //          .ready
		.in_data              (id_router_002_src_data),              //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_001_src_data),          //          .data
		.out_channel          (width_adapter_001_src_channel),       //          .channel
		.out_valid            (width_adapter_001_src_valid),         //          .valid
		.out_ready            (width_adapter_001_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (60),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (69),
		.IN_PKT_BYTE_CNT_L             (67),
		.IN_PKT_TRANS_COMPRESSED_READ  (61),
		.IN_PKT_BURSTWRAP_H            (72),
		.IN_PKT_BURSTWRAP_L            (70),
		.IN_PKT_BURST_SIZE_H           (75),
		.IN_PKT_BURST_SIZE_L           (73),
		.IN_PKT_RESPONSE_STATUS_H      (101),
		.IN_PKT_RESPONSE_STATUS_L      (100),
		.IN_PKT_TRANS_EXCLUSIVE        (66),
		.IN_PKT_BURST_TYPE_H           (77),
		.IN_PKT_BURST_TYPE_L           (76),
		.IN_ST_DATA_W                  (102),
		.OUT_PKT_ADDR_H                (42),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (51),
		.OUT_PKT_BYTE_CNT_L            (49),
		.OUT_PKT_TRANS_COMPRESSED_READ (43),
		.OUT_PKT_BURST_SIZE_H          (57),
		.OUT_PKT_BURST_SIZE_L          (55),
		.OUT_PKT_RESPONSE_STATUS_H     (83),
		.OUT_PKT_RESPONSE_STATUS_L     (82),
		.OUT_PKT_TRANS_EXCLUSIVE       (48),
		.OUT_PKT_BURST_TYPE_H          (59),
		.OUT_PKT_BURST_TYPE_L          (58),
		.OUT_ST_DATA_W                 (84),
		.ST_CHANNEL_W                  (20),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_002 (
		.clk                  (altpll_0_c1_clk),                     //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (cmd_xbar_mux_003_src_valid),          //      sink.valid
		.in_channel           (cmd_xbar_mux_003_src_channel),        //          .channel
		.in_startofpacket     (cmd_xbar_mux_003_src_startofpacket),  //          .startofpacket
		.in_endofpacket       (cmd_xbar_mux_003_src_endofpacket),    //          .endofpacket
		.in_ready             (cmd_xbar_mux_003_src_ready),          //          .ready
		.in_data              (cmd_xbar_mux_003_src_data),           //          .data
		.out_endofpacket      (width_adapter_002_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_002_src_data),          //          .data
		.out_channel          (width_adapter_002_src_channel),       //          .channel
		.out_valid            (width_adapter_002_src_valid),         //          .valid
		.out_ready            (width_adapter_002_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_002_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (42),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (51),
		.IN_PKT_BYTE_CNT_L             (49),
		.IN_PKT_TRANS_COMPRESSED_READ  (43),
		.IN_PKT_BURSTWRAP_H            (54),
		.IN_PKT_BURSTWRAP_L            (52),
		.IN_PKT_BURST_SIZE_H           (57),
		.IN_PKT_BURST_SIZE_L           (55),
		.IN_PKT_RESPONSE_STATUS_H      (83),
		.IN_PKT_RESPONSE_STATUS_L      (82),
		.IN_PKT_TRANS_EXCLUSIVE        (48),
		.IN_PKT_BURST_TYPE_H           (59),
		.IN_PKT_BURST_TYPE_L           (58),
		.IN_ST_DATA_W                  (84),
		.OUT_PKT_ADDR_H                (60),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (69),
		.OUT_PKT_BYTE_CNT_L            (67),
		.OUT_PKT_TRANS_COMPRESSED_READ (61),
		.OUT_PKT_BURST_SIZE_H          (75),
		.OUT_PKT_BURST_SIZE_L          (73),
		.OUT_PKT_RESPONSE_STATUS_H     (101),
		.OUT_PKT_RESPONSE_STATUS_L     (100),
		.OUT_PKT_TRANS_EXCLUSIVE       (66),
		.OUT_PKT_BURST_TYPE_H          (77),
		.OUT_PKT_BURST_TYPE_L          (76),
		.OUT_ST_DATA_W                 (102),
		.ST_CHANNEL_W                  (20),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_003 (
		.clk                  (altpll_0_c1_clk),                     //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (id_router_003_src_valid),             //      sink.valid
		.in_channel           (id_router_003_src_channel),           //          .channel
		.in_startofpacket     (id_router_003_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_003_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_003_src_ready),             //          .ready
		.in_data              (id_router_003_src_data),              //          .data
		.out_endofpacket      (width_adapter_003_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_003_src_data),          //          .data
		.out_channel          (width_adapter_003_src_channel),       //          .channel
		.out_valid            (width_adapter_003_src_valid),         //          .valid
		.out_ready            (width_adapter_003_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_003_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (60),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (69),
		.IN_PKT_BYTE_CNT_L             (67),
		.IN_PKT_TRANS_COMPRESSED_READ  (61),
		.IN_PKT_BURSTWRAP_H            (72),
		.IN_PKT_BURSTWRAP_L            (70),
		.IN_PKT_BURST_SIZE_H           (75),
		.IN_PKT_BURST_SIZE_L           (73),
		.IN_PKT_RESPONSE_STATUS_H      (101),
		.IN_PKT_RESPONSE_STATUS_L      (100),
		.IN_PKT_TRANS_EXCLUSIVE        (66),
		.IN_PKT_BURST_TYPE_H           (77),
		.IN_PKT_BURST_TYPE_L           (76),
		.IN_ST_DATA_W                  (102),
		.OUT_PKT_ADDR_H                (33),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (42),
		.OUT_PKT_BYTE_CNT_L            (40),
		.OUT_PKT_TRANS_COMPRESSED_READ (34),
		.OUT_PKT_BURST_SIZE_H          (48),
		.OUT_PKT_BURST_SIZE_L          (46),
		.OUT_PKT_RESPONSE_STATUS_H     (74),
		.OUT_PKT_RESPONSE_STATUS_L     (73),
		.OUT_PKT_TRANS_EXCLUSIVE       (39),
		.OUT_PKT_BURST_TYPE_H          (50),
		.OUT_PKT_BURST_TYPE_L          (49),
		.OUT_ST_DATA_W                 (75),
		.ST_CHANNEL_W                  (20),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_004 (
		.clk                  (altpll_0_c1_clk),                     //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (cmd_xbar_mux_005_src_valid),          //      sink.valid
		.in_channel           (cmd_xbar_mux_005_src_channel),        //          .channel
		.in_startofpacket     (cmd_xbar_mux_005_src_startofpacket),  //          .startofpacket
		.in_endofpacket       (cmd_xbar_mux_005_src_endofpacket),    //          .endofpacket
		.in_ready             (cmd_xbar_mux_005_src_ready),          //          .ready
		.in_data              (cmd_xbar_mux_005_src_data),           //          .data
		.out_endofpacket      (width_adapter_004_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_004_src_data),          //          .data
		.out_channel          (width_adapter_004_src_channel),       //          .channel
		.out_valid            (width_adapter_004_src_valid),         //          .valid
		.out_ready            (width_adapter_004_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_004_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (33),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (42),
		.IN_PKT_BYTE_CNT_L             (40),
		.IN_PKT_TRANS_COMPRESSED_READ  (34),
		.IN_PKT_BURSTWRAP_H            (45),
		.IN_PKT_BURSTWRAP_L            (43),
		.IN_PKT_BURST_SIZE_H           (48),
		.IN_PKT_BURST_SIZE_L           (46),
		.IN_PKT_RESPONSE_STATUS_H      (74),
		.IN_PKT_RESPONSE_STATUS_L      (73),
		.IN_PKT_TRANS_EXCLUSIVE        (39),
		.IN_PKT_BURST_TYPE_H           (50),
		.IN_PKT_BURST_TYPE_L           (49),
		.IN_ST_DATA_W                  (75),
		.OUT_PKT_ADDR_H                (60),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (69),
		.OUT_PKT_BYTE_CNT_L            (67),
		.OUT_PKT_TRANS_COMPRESSED_READ (61),
		.OUT_PKT_BURST_SIZE_H          (75),
		.OUT_PKT_BURST_SIZE_L          (73),
		.OUT_PKT_RESPONSE_STATUS_H     (101),
		.OUT_PKT_RESPONSE_STATUS_L     (100),
		.OUT_PKT_TRANS_EXCLUSIVE       (66),
		.OUT_PKT_BURST_TYPE_H          (77),
		.OUT_PKT_BURST_TYPE_L          (76),
		.OUT_ST_DATA_W                 (102),
		.ST_CHANNEL_W                  (20),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_005 (
		.clk                  (altpll_0_c1_clk),                     //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (id_router_005_src_valid),             //      sink.valid
		.in_channel           (id_router_005_src_channel),           //          .channel
		.in_startofpacket     (id_router_005_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_005_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_005_src_ready),             //          .ready
		.in_data              (id_router_005_src_data),              //          .data
		.out_endofpacket      (width_adapter_005_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_005_src_data),          //          .data
		.out_channel          (width_adapter_005_src_channel),       //          .channel
		.out_valid            (width_adapter_005_src_valid),         //          .valid
		.out_ready            (width_adapter_005_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_005_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (60),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (69),
		.IN_PKT_BYTE_CNT_L             (67),
		.IN_PKT_TRANS_COMPRESSED_READ  (61),
		.IN_PKT_BURSTWRAP_H            (72),
		.IN_PKT_BURSTWRAP_L            (70),
		.IN_PKT_BURST_SIZE_H           (75),
		.IN_PKT_BURST_SIZE_L           (73),
		.IN_PKT_RESPONSE_STATUS_H      (101),
		.IN_PKT_RESPONSE_STATUS_L      (100),
		.IN_PKT_TRANS_EXCLUSIVE        (66),
		.IN_PKT_BURST_TYPE_H           (77),
		.IN_PKT_BURST_TYPE_L           (76),
		.IN_ST_DATA_W                  (102),
		.OUT_PKT_ADDR_H                (33),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (42),
		.OUT_PKT_BYTE_CNT_L            (40),
		.OUT_PKT_TRANS_COMPRESSED_READ (34),
		.OUT_PKT_BURST_SIZE_H          (48),
		.OUT_PKT_BURST_SIZE_L          (46),
		.OUT_PKT_RESPONSE_STATUS_H     (74),
		.OUT_PKT_RESPONSE_STATUS_L     (73),
		.OUT_PKT_TRANS_EXCLUSIVE       (39),
		.OUT_PKT_BURST_TYPE_H          (50),
		.OUT_PKT_BURST_TYPE_L          (49),
		.OUT_ST_DATA_W                 (75),
		.ST_CHANNEL_W                  (20),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_006 (
		.clk                  (altpll_0_c1_clk),                        //       clk.clk
		.reset                (rst_controller_reset_out_reset),         // clk_reset.reset
		.in_valid             (cmd_xbar_demux_001_src10_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_001_src10_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_001_src10_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_001_src10_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_001_src10_ready),         //          .ready
		.in_data              (cmd_xbar_demux_001_src10_data),          //          .data
		.out_endofpacket      (width_adapter_006_src_endofpacket),      //       src.endofpacket
		.out_data             (width_adapter_006_src_data),             //          .data
		.out_channel          (width_adapter_006_src_channel),          //          .channel
		.out_valid            (width_adapter_006_src_valid),            //          .valid
		.out_ready            (width_adapter_006_src_ready),            //          .ready
		.out_startofpacket    (width_adapter_006_src_startofpacket),    //          .startofpacket
		.in_command_size_data (3'b000)                                  // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (33),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (42),
		.IN_PKT_BYTE_CNT_L             (40),
		.IN_PKT_TRANS_COMPRESSED_READ  (34),
		.IN_PKT_BURSTWRAP_H            (45),
		.IN_PKT_BURSTWRAP_L            (43),
		.IN_PKT_BURST_SIZE_H           (48),
		.IN_PKT_BURST_SIZE_L           (46),
		.IN_PKT_RESPONSE_STATUS_H      (74),
		.IN_PKT_RESPONSE_STATUS_L      (73),
		.IN_PKT_TRANS_EXCLUSIVE        (39),
		.IN_PKT_BURST_TYPE_H           (50),
		.IN_PKT_BURST_TYPE_L           (49),
		.IN_ST_DATA_W                  (75),
		.OUT_PKT_ADDR_H                (60),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (69),
		.OUT_PKT_BYTE_CNT_L            (67),
		.OUT_PKT_TRANS_COMPRESSED_READ (61),
		.OUT_PKT_BURST_SIZE_H          (75),
		.OUT_PKT_BURST_SIZE_L          (73),
		.OUT_PKT_RESPONSE_STATUS_H     (101),
		.OUT_PKT_RESPONSE_STATUS_L     (100),
		.OUT_PKT_TRANS_EXCLUSIVE       (66),
		.OUT_PKT_BURST_TYPE_H          (77),
		.OUT_PKT_BURST_TYPE_L          (76),
		.OUT_ST_DATA_W                 (102),
		.ST_CHANNEL_W                  (20),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_007 (
		.clk                  (altpll_0_c1_clk),                     //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (id_router_010_src_valid),             //      sink.valid
		.in_channel           (id_router_010_src_channel),           //          .channel
		.in_startofpacket     (id_router_010_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_010_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_010_src_ready),             //          .ready
		.in_data              (id_router_010_src_data),              //          .data
		.out_endofpacket      (width_adapter_007_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_007_src_data),          //          .data
		.out_channel          (width_adapter_007_src_channel),       //          .channel
		.out_valid            (width_adapter_007_src_valid),         //          .valid
		.out_ready            (width_adapter_007_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_007_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (102),
		.BITS_PER_SYMBOL     (102),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (20),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser (
		.in_clk            (altpll_0_c1_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (clk_clk),                               //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src6_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src6_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src6_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src6_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src6_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src6_data),          //              .data
		.out_ready         (crosser_out_ready),                     //           out.ready
		.out_valid         (crosser_out_valid),                     //              .valid
		.out_startofpacket (crosser_out_startofpacket),             //              .startofpacket
		.out_endofpacket   (crosser_out_endofpacket),               //              .endofpacket
		.out_channel       (crosser_out_channel),                   //              .channel
		.out_data          (crosser_out_data),                      //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (102),
		.BITS_PER_SYMBOL     (102),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (20),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_001 (
		.in_clk            (altpll_0_c1_clk),                        //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),         //  in_clk_reset.reset
		.out_clk           (up_clocks_1_audio_clk_clk),              //       out_clk.clk
		.out_reset         (rst_controller_002_reset_out_reset),     // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src13_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src13_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src13_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src13_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src13_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src13_data),          //              .data
		.out_ready         (crosser_001_out_ready),                  //           out.ready
		.out_valid         (crosser_001_out_valid),                  //              .valid
		.out_startofpacket (crosser_001_out_startofpacket),          //              .startofpacket
		.out_endofpacket   (crosser_001_out_endofpacket),            //              .endofpacket
		.out_channel       (crosser_001_out_channel),                //              .channel
		.out_data          (crosser_001_out_data),                   //              .data
		.in_empty          (1'b0),                                   //   (terminated)
		.in_error          (1'b0),                                   //   (terminated)
		.out_empty         (),                                       //   (terminated)
		.out_error         ()                                        //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (102),
		.BITS_PER_SYMBOL     (102),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (20),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_002 (
		.in_clk            (altpll_0_c1_clk),                        //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),         //  in_clk_reset.reset
		.out_clk           (up_clocks_1_audio_clk_clk),              //       out_clk.clk
		.out_reset         (rst_controller_002_reset_out_reset),     // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src14_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src14_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src14_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src14_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src14_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src14_data),          //              .data
		.out_ready         (crosser_002_out_ready),                  //           out.ready
		.out_valid         (crosser_002_out_valid),                  //              .valid
		.out_startofpacket (crosser_002_out_startofpacket),          //              .startofpacket
		.out_endofpacket   (crosser_002_out_endofpacket),            //              .endofpacket
		.out_channel       (crosser_002_out_channel),                //              .channel
		.out_data          (crosser_002_out_data),                   //              .data
		.in_empty          (1'b0),                                   //   (terminated)
		.in_error          (1'b0),                                   //   (terminated)
		.out_empty         (),                                       //   (terminated)
		.out_error         ()                                        //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (102),
		.BITS_PER_SYMBOL     (102),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (20),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_003 (
		.in_clk            (clk_clk),                               //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (altpll_0_c1_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_006_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_006_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_006_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_006_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_006_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_006_src0_data),          //              .data
		.out_ready         (crosser_003_out_ready),                 //           out.ready
		.out_valid         (crosser_003_out_valid),                 //              .valid
		.out_startofpacket (crosser_003_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_003_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_003_out_channel),               //              .channel
		.out_data          (crosser_003_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (102),
		.BITS_PER_SYMBOL     (102),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (20),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_004 (
		.in_clk            (up_clocks_1_audio_clk_clk),             //        in_clk.clk
		.in_reset          (rst_controller_002_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (altpll_0_c1_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_013_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_013_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_013_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_013_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_013_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_013_src0_data),          //              .data
		.out_ready         (crosser_004_out_ready),                 //           out.ready
		.out_valid         (crosser_004_out_valid),                 //              .valid
		.out_startofpacket (crosser_004_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_004_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_004_out_channel),               //              .channel
		.out_data          (crosser_004_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (102),
		.BITS_PER_SYMBOL     (102),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (20),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_005 (
		.in_clk            (up_clocks_1_audio_clk_clk),             //        in_clk.clk
		.in_reset          (rst_controller_002_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (altpll_0_c1_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_014_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_014_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_014_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_014_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_014_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_014_src0_data),          //              .data
		.out_ready         (crosser_005_out_ready),                 //           out.ready
		.out_valid         (crosser_005_out_valid),                 //              .valid
		.out_startofpacket (crosser_005_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_005_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_005_out_channel),               //              .channel
		.out_data          (crosser_005_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	niosII_system_irq_mapper irq_mapper (
		.clk           (altpll_0_c1_clk),                //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (nios2_qsys_0_d_irq_irq)          //    sender.irq
	);

endmodule
